library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity fsub_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity fsub_tb;

architecture testbench of fsub_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "00111111100000000000000000000000",
    1 => "00111111011100001000111111111101",
    2 => "00111110101100101011011111111111",
    3 => "00111110101011110001110010010000",
    4 => "00111111100000000000000000000000",
    5 => "00111111010111011011010111111010",
    6 => "00111111000001100000100111111111",
    7 => "00111110111111111111111101000111",
    8 => "00000000000000000000000000000000",
    9 => "00000000000000000000000000000000",
    10 => "00000000000000000000000000000000",
    11 => "11000010100011000000000000000000",
    12 => "01000010000011000000000000000000",
    13 => "11000001101000000000000000000000",
    14 => "00111111110010010000111111011000",
    15 => "00111111100000000000000000000000",
    16 => "00111111010001000010010101001010",
    17 => "00000000000000000000000000000000",
    18 => "00111111110010010000111111011000",
    19 => "00111111001100101011100110110010",
    20 => "00111111001001001000111101111010",
    21 => "00111111110010010000111111011000",
    22 => "00111111100000000000000000000000",
    23 => "00111111010001000010010101001010",
    24 => "00111111110010010000111111011000",
    25 => "00111111001100101011100110110010",
    26 => "00111111001001001000111101111010",
    27 => "00000000000000000000000000000000",
    28 => "00000000000000000000000000000000",
    29 => "00111111111001100110011001100111",
    30 => "00111101110000000010001000111101",
    31 => "10111110000100110001011000100111",
    32 => "00111111101010010111100010100100",
    33 => "10111110000001100000101011000010",
    34 => "10111110000001011010100011011000",
    35 => "00000000000000000000000000000000",
    36 => "00111111100000000000000000000000",
    37 => "00111111011111011100111101010011",
    38 => "00000000000000000000000000000000",
    39 => "00111101101111100111110101101111",
    40 => "10111110000101000110011110101011",
    41 => "00111111101010000010011010100001",
    42 => "00111111110010010000111111011000",
    43 => "00111111100000000000000000000000",
    44 => "00111111011010111001100001111101",
    45 => "00111111110010010000111111011000",
    46 => "00111110110011011100111111001000",
    47 => "00111110110010000101000001010010",
    48 => "00111101000101010011111110011000",
    49 => "10111110000000010100101010110010",
    50 => "00111111011011000101100000010001",
    51 => "10111101101110100000000101011000",
    52 => "10111101101110011011111111101000",
    53 => "00000000000000000000000000000000",
    54 => "00111111100000000000000000000000",
    55 => "00111111011111101111000111100100",
    56 => "00000000000000000000000000000000",
    57 => "00111101101110110000111101011000",
    58 => "10111110000101110000001101001011",
    59 => "00111111101001011010010110001001",
    60 => "00111111110010010000111111011000",
    61 => "00111111100000000000000000000000",
    62 => "00111111011010011100101111001100",
    63 => "00111111110010010000111111011000",
    64 => "00111110110101101101001110111000",
    65 => "00111110110100001001010000111111",
    66 => "00111101000110010001001010010111",
    67 => "10111110000000110110011001111010",
    68 => "00111111011100000001101010111101",
    69 => "10111101101111010000001101111011",
    70 => "10111101101111001011111011010001",
    71 => "00000000000000000000000000000000",
    72 => "00111111100000000000000000000000",
    73 => "00111111011111101110100100010110",
    74 => "00000000000000000000000000000000",
    75 => "00111101101110110010011000001000",
    76 => "10111110000101101111001010101011",
    77 => "00111111101001011011010100001110",
    78 => "00111111110010010000111111011000",
    79 => "00111111100000000000000000000000",
    80 => "00111111011010011101011100101011",
    81 => "00111111110010010000111111011000",
    82 => "00111110110101101001101111011100",
    83 => "00111110110100000110000100111010",
    84 => "00111101000110001111110001101110",
    85 => "10111110000000110101101001101110",
    86 => "00111111011100000000010101010010",
    87 => "10111101101111001111001001011001",
    88 => "10111101101111001010110111000001",
    89 => "00000000000000000000000000000000",
    90 => "00111111100000000000000000000000",
    91 => "00111111011111101110100101001000",
    92 => "00000000000000000000000000000000",
    93 => "00111101101110110010010110000011",
    94 => "10111110000101101111001100001100",
    95 => "00111111101001011011010010110110",
    96 => "00111111110010010000111111011000",
    97 => "00111111100000000000000000000000",
    98 => "00111111011010011101011011101011",
    99 => "00111111110010010000111111011000",
    100 => "00111110110101101001110100011000",
    101 => "00111110110100000110001001011010",
    102 => "00111101000110001111110011101011",
    103 => "10111110000000110101101010110010",
    104 => "00111111011100000000010111001100",
    105 => "10111101101111001111001010111011",
    106 => "10111101101111001010111000100011",
    107 => "00000000000000000000000000000000",
    108 => "00111111100000000000000000000000",
    109 => "00111111011111101110100101001000",
    110 => "00000000000000000000000000000000",
    111 => "00111101101110110010010110000111",
    112 => "10111110000101101111001100001001",
    113 => "00111111101001011011010010110111",
    114 => "00111111110010010000111111011000",
    115 => "00111111100000000000000000000000",
    116 => "00111111011010011101011011101011",
    117 => "00111111110010010000111111011000",
    118 => "00111110110101101001110100010100",
    119 => "00111110110100000110001001010111",
    120 => "00000000000000000000000000000000",
    121 => "00000000000000000000000000000000",
    122 => "00000000000000000000000000000000",
    123 => "00111101110000000010001000111101",
    124 => "10111110000100110001011000100111",
    125 => "00111111101010010111100010100100",
    126 => "00111111110010010000111111011000",
    127 => "00111111100000000000000000000000",
    128 => "00111111011011001000001111011110",
    129 => "00111111110010010000111111011000",
    130 => "00111110110010010000111011111000",
    131 => "00111110110000111110111001001101",
    132 => "00111101000100110000110011100101",
    133 => "10111110000000000000110101111001",
    134 => "00111111011010100001111101011011",
    135 => "00111111110010010000111111011000",
    136 => "00111111100000000000000000000000",
    137 => "00111111001110010110101000011001",
    138 => "00111111110010010000111111011000",
    139 => "00111111010000101101111000000011",
    140 => "00111111001100001001100000000110",
    141 => "00111101000000111010000000001001",
    142 => "10111101111011011001100000111101",
    143 => "00111111010110010100101111001111",
    144 => "00111111010000000001110011100001",
    145 => "00111111001011101001011010111000",
    146 => "00111111100000000000000000000000",
    147 => "00111111001110110100110001010000",
    148 => "00111101000001001000000110111011",
    149 => "10111101111011101011010010010011",
    150 => "00111111010110100101000011101001",
    151 => "00111111010000010000011111100000",
    152 => "00111111001011110100001001011100",
    153 => "00111111100000000000000000000000",
    154 => "00111111001110101010110000110110",
    155 => "00111101000001000111001001110101",
    156 => "10111101111011101010000101100100",
    157 => "00111111010110100011111101001100",
    158 => "00111111010000001111100000000101",
    159 => "00111111001011110011011011001101",
    160 => "00111111100000000000000000000000",
    161 => "00111111001110101011011100001000",
    162 => "00111101000001000111001101110111",
    163 => "10111101111011101010001010101000",
    164 => "00111111010110100100000001110110",
    165 => "00111111010000001111100100010011",
    166 => "00111111001011110011011110010001",
    167 => "00111111100000000000000000000000",
    168 => "00111111001110101011011001001111",
    169 => "00111101000001000111001101100110",
    170 => "10111101111011101010001010010011",
    171 => "00111111010110100100000001100011",
    172 => "00111111010000001111100100000000",
    173 => "00111111001011110011011110000011",
    174 => "00111111100000000000000000000000",
    175 => "00111111001110101011011001011100",
    176 => "00111101000001000111001101101000",
    177 => "10111101111011101010001010010101",
    178 => "00111111010110100100000001100101",
    179 => "00111111010000001111100100000011",
    180 => "00111111001011110011011110000110",
    181 => "00111111100000000000000000000000",
    182 => "00111111001110101011011001011010",
    183 => "00111101000001000111001101100110",
    184 => "10111101111011101010001010010011",
    185 => "00111111010110100100000001100011",
    186 => "00111111010000001111100100000000",
    187 => "00111111001011110011011110000011",
    188 => "00111111100000000000000000000000",
    189 => "00111111001110101011011001011100",
    190 => "00111101000001000111001101101000",
    191 => "10111101111011101010001010010101",
    192 => "00111111010110100100000001100101",
    193 => "00111111010000001111100100000011",
    194 => "00111111001011110011011110000110",
    195 => "00111111100000000000000000000000",
    196 => "00111111001110101011011001011010",
    197 => "00000000000000000000000000000000",
    198 => "00000000000000000000000000000000",
    199 => "00000000000000000000000000000000",
    200 => "00111111000110011001100110011010",
    201 => "00111101110000000010001000111101",
    202 => "10111110000100110001011000100111",
    203 => "00111111101010010111100010100100",
    204 => "10111110110010010001000000100010",
    205 => "10111110110000111110111101011111",
    206 => "00000000000000000000000000000000",
    207 => "00111111100000000000000000000000",
    208 => "00111111011011001000001110100101",
    209 => "00000000000000000000000000000000",
    210 => "00111101101100011000001000011111",
    211 => "10111110000111010100000100110101",
    212 => "00111111101000000011101000101000",
    213 => "00111111110010010000111111011000",
    214 => "00111111100000000000000000000000",
    215 => "00111111011001011010011110010110",
    216 => "00111111110010010000111111011000",
    217 => "00111110111010100101011001001100",
    218 => "00111110111000100011110111000100",
    219 => "00111101000111110010101001101000",
    220 => "10111110000001101010001010101110",
    221 => "00111111011101011101001010001111",
    222 => "10111110100100010011000011100110",
    223 => "10111110100011110100000010111110",
    224 => "00000000000000000000000000000000",
    225 => "00111111100000000000000000000000",
    226 => "00111111011101011100011010011010",
    227 => "00000000000000000000000000000000",
    228 => "00111101100111010010001011111111",
    229 => "10111110001001011000110011111110",
    230 => "00111111100110011110001111010110",
    231 => "00111111110010010000111111011000",
    232 => "00111111100000000000000000000000",
    233 => "00111111011000000110001111101011",
    234 => "00111111110010010000111111011000",
    235 => "00111111000000001001001101010010",
    236 => "00111110111101100111100111100001",
    237 => "00111101000111010111001110101101",
    238 => "10111110000001011011110110101111",
    239 => "00111111011101000011111101111110",
    240 => "10111110100100000011111100001111",
    241 => "10111110100011100101100001111111",
    242 => "00000000000000000000000000000000",
    243 => "00111111100000000000000000000000",
    244 => "00111111011101011110100001010100",
    245 => "00000000000000000000000000000000",
    246 => "00111101100111001110111001110011",
    247 => "10111110001001011001100101111110",
    248 => "00111111100110011101100100101110",
    249 => "00111111110010010000111111011000",
    250 => "00111111100000000000000000000000",
    251 => "00111111011000000101101010110000",
    252 => "00111111110010010000111111011000",
    253 => "00111111000000001010011010000000",
    254 => "00111110111101101001101110000000",
    255 => "00111101000111010101111100010110",
    256 => "10111110000001011011001011011100",
    257 => "00111111011101000010110001101001",
    258 => "10111110100100000011001110011011",
    259 => "10111110100011100100110110000000",
    260 => "00000000000000000000000000000000",
    261 => "00111111100000000000000000000000",
    262 => "00111111011101011110100111101011",
    263 => "00000000000000000000000000000000",
    264 => "00111101100111001110101111111101",
    265 => "10111110001001011001101000010010",
    266 => "00111111100110011101100010101111",
    267 => "00111111110010010000111111011000",
    268 => "00111111100000000000000000000000",
    269 => "00111111011000000101101001000001",
    270 => "00111111110010010000111111011000",
    271 => "00111111000000001010011101100110",
    272 => "00111110111101101001110100010011",
    273 => "00111101000111010101111000100000",
    274 => "10111110000001011011001001011010",
    275 => "00111111011101000010101110000101",
    276 => "10111110100100000011001100010011",
    277 => "10111110100011100100110011111100",
    278 => "00000000000000000000000000000000",
    279 => "00111111100000000000000000000000",
    280 => "00111111011101011110100111111110",
    281 => "00000000000000000000000000000000",
    282 => "00111101100111001110101111100000",
    283 => "10111110001001011001101000011001",
    284 => "00111111100110011101100010101001",
    285 => "00111111110010010000111111011000",
    286 => "00111111100000000000000000000000",
    287 => "00111111011000000101101000111100",
    288 => "00111111110010010000111111011000",
    289 => "00111111000000001010011101110000",
    290 => "00111110111101101001110100100100",
    291 => "00000000000000000000000000000000",
    292 => "00000000000000000000000000000000",
    293 => "00000000000000000000000000000000",
    294 => "00111101110000000010001000111101",
    295 => "10111110000100110001011000100111",
    296 => "00111111101010010111100010100100",
    297 => "00111111110010010000111111011000",
    298 => "00111111100000000000000000000000",
    299 => "00111111010010110010000001111101",
    300 => "00111111110010010000111111011000",
    301 => "00111111001001111000110011011011",
    302 => "00111111000110111101100000101010",
    303 => "00111101011010011110110011110000",
    304 => "10111110001000011110010011101110",
    305 => "00111111100100010110111001011101",
    306 => "00111111110010010000111111011000",
    307 => "00111111100000000000000000000000",
    308 => "00111111010110001010110001101100",
    309 => "00111111110010010000111111011000",
    310 => "00111111000011111100110100101100",
    311 => "00111111000010000101101110111110",
    312 => "00111101000010010111101001000110",
    313 => "10111101111101001101100100101010",
    314 => "00111111010111111110111101010111",
    315 => "00111111000110100001000101111000",
    316 => "00111111000100001110111110100100",
    317 => "00111111100000000000000000000000",
    318 => "00111111010100110000100110110010",
    319 => "00111101001100011000011000001000",
    320 => "10111110000011110111010110010100",
    321 => "00111111100000101000011001100101",
    322 => "00111111110010010000111111011000",
    323 => "00111111100000000000000000000000",
    324 => "00111111010010010011110100110100",
    325 => "00111111110010010000111111011000",
    326 => "00111111001010101010000111101010",
    327 => "00111111000111100100011101011010",
    328 => "00111101000000110011111100111000",
    329 => "10111101111011010001110111000010",
    330 => "00111111010110001101101100111110",
    331 => "00111111000101010001110100000001",
    332 => "00111111000011001101001100010110",
    333 => "00111111100000000000000000000000",
    334 => "00111111010101011100110011101001",
    335 => "00111101001100001110001001001010",
    336 => "10111110000011110010110011011001",
    337 => "00111111100000100100100011010101",
    338 => "00111111110010010000111111011000",
    339 => "00111111100000000000000000000000",
    340 => "00111111010010001111100010111100",
    341 => "00111111110010010000111111011000",
    342 => "00111111001010110001000010111011",
    343 => "00111111000111101001111001101000",
    344 => "00111101000000110011101101010011",
    345 => "10111101111011010001100011010011",
    346 => "00111111010110001101011010110101",
    347 => "00111111000101010001100111010100",
    348 => "00111111000011001101000001101110",
    349 => "00111111100000000000000000000000",
    350 => "00111111010101011100111010101000",
    351 => "00111101001100001110000111101111",
    352 => "10111110000011110010110010110000",
    353 => "00111111100000100100100010110100",
    354 => "00111111110010010000111111011000",
    355 => "00111111100000000000000000000000",
    356 => "00111111010010001111100010011000",
    357 => "00111111110010010000111111011000",
    358 => "00111111001010110001000011110110",
    359 => "00111111000111101001111010010110",
    360 => "00111101000000110011101101001111",
    361 => "10111101111011010001100011001110",
    362 => "00111111010110001101011010110001",
    363 => "00111111000101010001100111010001",
    364 => "00111111000011001101000001101100",
    365 => "00111111100000000000000000000000",
    366 => "00111111010101011100111010101010",
    367 => "00111101001100001110000111101010",
    368 => "10111110000011110010110010101101",
    369 => "00111111100000100100100010110010",
    370 => "00111111110010010000111111011000",
    371 => "00111111100000000000000000000000",
    372 => "00111111010010001111100010010101",
    373 => "00111111110010010000111111011000",
    374 => "00111111001010110001000011111010",
    375 => "00111111000111101001111010011001",
    376 => "00000000000000000000000000000000",
    377 => "00000000000000000000000000000000",
    378 => "00000000000000000000000000000000",
    379 => "00111110110011001100110011001110",
    380 => "00111101110000000010001000111101",
    381 => "10111110000100110001011000100111",
    382 => "00111111101010010111100010100100",
    383 => "10111111001001111000110101110001",
    384 => "10111111000110111101100010100001",
    385 => "00000000000000000000000000000000",
    386 => "00111111100000000000000000000000",
    387 => "00111111010010110010000000100010",
    388 => "00000000000000000000000000000000",
    389 => "00111101100110000110110111111000",
    390 => "10111110001001100111111100000110",
    391 => "00111111100110001111111001100101",
    392 => "00111111110010010000111111011000",
    393 => "00111111100000000000000000000000",
    394 => "00111111010111111001110000010100",
    395 => "00111111110010010000111111011000",
    396 => "00111111000000100011000001010010",
    397 => "00111110111110010100110010100010",
    398 => "00111101000110110110110010010000",
    399 => "10111110000001001010101010111100",
    400 => "00111111011100100101100111010100",
    401 => "10111110111011101000001101110000",
    402 => "10111110111001011111101011110010",
    403 => "00000000000000000000000000000000",
    404 => "00111111100000000000000000000000",
    405 => "00111111011001001011100110000010",
    406 => "00000000000000000000000000000000",
    407 => "00111101011100001101111101001111",
    408 => "10111110001000110100001001101001",
    409 => "00111111100100101000100001001101",
    410 => "00111111110010010000111111011000",
    411 => "00111111100000000000000000000000",
    412 => "00111111010110011011100011010111",
    413 => "00111111110010010000111111011000",
    414 => "00111111000011011101000110110000",
    415 => "00111111000001101010110100101100",
    416 => "00111101000010101110110010010101",
    417 => "10111101111101101001100100000011",
    418 => "00111111011000011000011100100001",
    419 => "10111110110111011011000010111100",
    420 => "10111110110101101101010000000110",
    421 => "00000000000000000000000000000000",
    422 => "00111111100000000000000000000000",
    423 => "00111111011010000110000010100101",
    424 => "00000000000000000000000000000000",
    425 => "00111101011011001011110001000000",
    426 => "10111110001000100111100001101001",
    427 => "00111111100100011110010001100011",
    428 => "00111111110010010000111111011000",
    429 => "00111111100000000000000000000000",
    430 => "00111111010110010001110100110010",
    431 => "00111111110010010000111111011000",
    432 => "00111111000011101111100010111010",
    433 => "00111111000001111010011111000000",
    434 => "00111101000010100000101111100110",
    435 => "10111101111101011000100111001111",
    436 => "00111111011000001001000001001010",
    437 => "10111110110111001011100111100110",
    438 => "10111110110101011111001111011110",
    439 => "00000000000000000000000000000000",
    440 => "00111111100000000000000000000000",
    441 => "00111111011010001001010001001111",
    442 => "00000000000000000000000000000000",
    443 => "00111101011011001000100000101010",
    444 => "10111110001000100110111000000010",
    445 => "00111111100100011101110000001000",
    446 => "00111111110010010000111111011000",
    447 => "00111111100000000000000000000000",
    448 => "00111111010110010001010100111010",
    449 => "00111111110010010000111111011000",
    450 => "00111111000011110000011111000110",
    451 => "00111111000001111011010010000010",
    452 => "00111101000010100000000100100010",
    453 => "10111101111101010111110011000101",
    454 => "00111111011000001000010001101010",
    455 => "10111110110111001010111000000110",
    456 => "10111110110101011110100100010100",
    457 => "00000000000000000000000000000000",
    458 => "00111111100000000000000000000000",
    459 => "00111111011010001001011011001010",
    460 => "00000000000000000000000000000000",
    461 => "00111101011011001000010110101111",
    462 => "10111110001000100110110110000011",
    463 => "00111111100100011101101110100010",
    464 => "00111111110010010000111111011000",
    465 => "00111111100000000000000000000000",
    466 => "00111111010110010001010011011001",
    467 => "00111111110010010000111111011000",
    468 => "00111111000011110000100001111100",
    469 => "00111111000001111011010100011100",
    470 => "00000000000000000000000000000000",
    471 => "00000000000000000000000000000000",
    472 => "00000000000000000000000000000000",
    473 => "00111101110000000010001000111101",
    474 => "10111110000100110001011000100111",
    475 => "00111111101010010111100010100100",
    476 => "00111111001001111000110101110100",
    477 => "00111111000110111101100010100011",
    478 => "00111111100000000000000000000000",
    479 => "00111111010010110010000000100000",
    480 => "00111101100110000110110111111000",
    481 => "10111110001001100111111100000110",
    482 => "00111111100110001111111001100101",
    483 => "00111111110010010000111111011000",
    484 => "00111111100000000000000000000000",
    485 => "00111111010111111001110000010100",
    486 => "00111111110010010000111111011000",
    487 => "00111111000000100011000001010010",
    488 => "00111110111110010100110010100010",
    489 => "00111101000110110110110010010000",
    490 => "10111110000001001010101010111100",
    491 => "00111111011100100101100111010100",
    492 => "00111110111011101000001101110011",
    493 => "00111110111001011111101011110101",
    494 => "00111111100000000000000000000000",
    495 => "00111111011001001011100110000001",
    496 => "00111101011100001101111101001100",
    497 => "10111110001000110100001001101001",
    498 => "00111111100100101000100001001100",
    499 => "00111111110010010000111111011000",
    500 => "00111111100000000000000000000000",
    501 => "00111111010110011011100011010110",
    502 => "00111111110010010000111111011000",
    503 => "00111111000011011101000110110010",
    504 => "00111111000001101010110100101110",
    505 => "00111101000010101110110010010101",
    506 => "10111101111101101001100100000011",
    507 => "00111111011000011000011100100001",
    508 => "00111110110111011011000010111111",
    509 => "00111110110101101101010000001001",
    510 => "00111111100000000000000000000000",
    511 => "00111111011010000110000010100101",
    512 => "00111101011011001011110000111110",
    513 => "10111110001000100111100001101000",
    514 => "00111111100100011110010001100100",
    515 => "00111111110010010000111111011000",
    516 => "00111111100000000000000000000000",
    517 => "00111111010110010001110100110010",
    518 => "00111111110010010000111111011000",
    519 => "00111111000011101111100010111000",
    520 => "00111111000001111010011110111110",
    521 => "00111101000010100000101111100101",
    522 => "10111101111101011000100111001101",
    523 => "00111111011000001001000001001001",
    524 => "00111110110111001011100111100111",
    525 => "00111110110101011111001111100000",
    526 => "00111111100000000000000000000000",
    527 => "00111111011010001001010001001110",
    528 => "00111101011011001000100000100100",
    529 => "10111110001000100110111000000001",
    530 => "00111111100100011101110000000110",
    531 => "00111111110010010000111111011000",
    532 => "00111111100000000000000000000000",
    533 => "00111111010110010001010100111000",
    534 => "00111111110010010000111111011000",
    535 => "00111111000011110000011111001000",
    536 => "00111111000001111011010010000011",
    537 => "00111101000010100000000100100010",
    538 => "10111101111101010111110011000101",
    539 => "00111111011000001000010001101010",
    540 => "00111110110111001010111000001001",
    541 => "00111110110101011110100100010111",
    542 => "00111111100000000000000000000000",
    543 => "00111111011010001001011011001001",
    544 => "00111101011011001000010110101100",
    545 => "10111110001000100110110110000010",
    546 => "00111111100100011101101110100010",
    547 => "00111111110010010000111111011000",
    548 => "00111111100000000000000000000000",
    549 => "00111111010110010001010011011001",
    550 => "00111111110010010000111111011000",
    551 => "00111111000011110000100001111100",
    552 => "00111111000001111011010100011100",
    553 => "00000000000000000000000000000000",
    554 => "00000000000000000000000000000000",
    555 => "00000000000000000000000000000000",
    556 => "00111110010011001100110011001110",
    557 => "00111101110000000010001000111101",
    558 => "10111110000100110001011000100111",
    559 => "00111111101010010111100010100100",
    560 => "10111111011010101001001011010011",
    561 => "10111111010010110010000001011000",
    562 => "00000000000000000000000000000000",
    563 => "00111111100000000000000000000000",
    564 => "00111111000111000000110001111010",
    565 => "00000000000000000000000000000000",
    566 => "00111101011010011110110011010010",
    567 => "10111110001000011110010011100111",
    568 => "00111111100100010110111001011001",
    569 => "00111111110010010000111111011000",
    570 => "00111111100000000000000000000000",
    571 => "00111111010110001010110001101000",
    572 => "00111111110010010000111111011000",
    573 => "00111111000011111100110100110100",
    574 => "00111111000010000101101111000101",
    575 => "00111101000010010111101000111110",
    576 => "10111101111101001101100100100001",
    577 => "00111111010111111110111101010000",
    578 => "10111111000110100001000101110010",
    579 => "10111111000100001110111110100000",
    580 => "00000000000000000000000000000000",
    581 => "00111111100000000000000000000000",
    582 => "00111111010100110000100110110100",
    583 => "00000000000000000000000000000000",
    584 => "00111101001100011000011000000100",
    585 => "10111110000011110111010110010011",
    586 => "00111111100000101000011001100100",
    587 => "00111111110010010000111111011000",
    588 => "00111111100000000000000000000000",
    589 => "00111111010010010011110100110010",
    590 => "00111111110010010000111111011000",
    591 => "00111111001010101010000111101100",
    592 => "00111111000111100100011101011011",
    593 => "00111101000000110011111100111000",
    594 => "10111101111011010001110111000010",
    595 => "00111111010110001101101100111110",
    596 => "10111111000101010001110011111111",
    597 => "10111111000011001101001100010100",
    598 => "00000000000000000000000000000000",
    599 => "00111111100000000000000000000000",
    600 => "00111111010101011100110011101011",
    601 => "00000000000000000000000000000000",
    602 => "00111101001100001110001001001110",
    603 => "10111110000011110010110011011010",
    604 => "00111111100000100100100011010111",
    605 => "00111111110010010000111111011000",
    606 => "00111111100000000000000000000000",
    607 => "00111111010010001111100010111111",
    608 => "00111111110010010000111111011000",
    609 => "00111111001010110001000010110111",
    610 => "00111111000111101001111001100100",
    611 => "00111101000000110011101101010011",
    612 => "10111101111011010001100011010011",
    613 => "00111111010110001101011010110101",
    614 => "10111111000101010001100111010010",
    615 => "10111111000011001101000001101110",
    616 => "00000000000000000000000000000000",
    617 => "00111111100000000000000000000000",
    618 => "00111111010101011100111010101001",
    619 => "00000000000000000000000000000000",
    620 => "00111101001100001110000111101101",
    621 => "10111110000011110010110010110000",
    622 => "00111111100000100100100010110010",
    623 => "00111111110010010000111111011000",
    624 => "00111111100000000000000000000000",
    625 => "00111111010010001111100010010101",
    626 => "00111111110010010000111111011000",
    627 => "00111111001010110001000011111010",
    628 => "00111111000111101001111010011001",
    629 => "00111101000000110011101101010011",
    630 => "10111101111011010001100011010011",
    631 => "00111111010110001101011010110101",
    632 => "10111111000101010001100111010010",
    633 => "10111111000011001101000001101110",
    634 => "00000000000000000000000000000000",
    635 => "00111111100000000000000000000000",
    636 => "00111111010101011100111010101001",
    637 => "00000000000000000000000000000000",
    638 => "00111101001100001110000111101101",
    639 => "10111110000011110010110010110000",
    640 => "00111111100000100100100010110010",
    641 => "00111111110010010000111111011000",
    642 => "00111111100000000000000000000000",
    643 => "00111111010010001111100010010101",
    644 => "00111111110010010000111111011000",
    645 => "00111111001010110001000011111010",
    646 => "00111111000111101001111010011001",
    647 => "00000000000000000000000000000000",
    648 => "00000000000000000000000000000000",
    649 => "00000000000000000000000000000000",
    650 => "00111101110000000010001000111101",
    651 => "10111110000100110001011000100111",
    652 => "00111111101010010111100010100100",
    653 => "00111110110010010001000000100100",
    654 => "00111110110000111110111101100001",
    655 => "00111111100000000000000000000000",
    656 => "00111111011011001000001110100101",
    657 => "00111101101100011000001000011111",
    658 => "10111110000111010100000100110101",
    659 => "00111111101000000011101000101000",
    660 => "00111111110010010000111111011000",
    661 => "00111111100000000000000000000000",
    662 => "00111111011001011010011110010110",
    663 => "00111111110010010000111111011000",
    664 => "00111110111010100101011001001100",
    665 => "00111110111000100011110111000100",
    666 => "00111101000111110010101001101000",
    667 => "10111110000001101010001010101110",
    668 => "00111111011101011101001010001111",
    669 => "00111110100100010011000011101000",
    670 => "00111110100011110100000011000000",
    671 => "00111111100000000000000000000000",
    672 => "00111111011101011100011010011010",
    673 => "00111101100111010010001011111101",
    674 => "10111110001001011000110011111110",
    675 => "00111111100110011110001111010110",
    676 => "00111111110010010000111111011000",
    677 => "00111111100000000000000000000000",
    678 => "00111111011000000110001111101011",
    679 => "00111111110010010000111111011000",
    680 => "00111111000000001001001101010010",
    681 => "00111110111101100111100111100001",
    682 => "00111101000111010111001110101101",
    683 => "10111110000001011011110110101111",
    684 => "00111111011101000011111101111110",
    685 => "00111110100100000011111100010001",
    686 => "00111110100011100101100010000001",
    687 => "00111111100000000000000000000000",
    688 => "00111111011101011110100001010100",
    689 => "00111101100111001110111001110001",
    690 => "10111110001001011001100101111110",
    691 => "00111111100110011101100100101110",
    692 => "00111111110010010000111111011000",
    693 => "00111111100000000000000000000000",
    694 => "00111111011000000101101010110000",
    695 => "00111111110010010000111111011000",
    696 => "00111111000000001010011010000000",
    697 => "00111110111101101001101110000000",
    698 => "00111101000111010101111100010110",
    699 => "10111110000001011011001011011100",
    700 => "00111111011101000010110001101001",
    701 => "00111110100100000011001110011101",
    702 => "00111110100011100100110110000010",
    703 => "00111111100000000000000000000000",
    704 => "00111111011101011110100111101011",
    705 => "00111101100111001110101111111101",
    706 => "10111110001001011001101000010010",
    707 => "00111111100110011101100010101111",
    708 => "00111111110010010000111111011000",
    709 => "00111111100000000000000000000000",
    710 => "00111111011000000101101001000001",
    711 => "00111111110010010000111111011000",
    712 => "00111111000000001010011101100110",
    713 => "00111110111101101001110100010011",
    714 => "00111101000111010101111000100000",
    715 => "10111110000001011011001001011010",
    716 => "00111111011101000010101110000101",
    717 => "00111110100100000011001100010101",
    718 => "00111110100011100100110011111110",
    719 => "00111111100000000000000000000000",
    720 => "00111111011101011110100111111110",
    721 => "00111101100111001110101111011110",
    722 => "10111110001001011001101000011010",
    723 => "00111111100110011101100010101000",
    724 => "00111111110010010000111111011000",
    725 => "00111111100000000000000000000000",
    726 => "00111111011000000101101000111100",
    727 => "00111111110010010000111111011000",
    728 => "00111111000000001010011101110010",
    729 => "00111110111101101001110100100111",
    730 => "00000000000000000000000000000000",
    731 => "00000000000000000000000000000000",
    732 => "00000000000000000000000000000000",
    733 => "00000000000000000000000000000000",
    734 => "00111101110000000010001000111101",
    735 => "10111110000100110001011000100111",
    736 => "00111111101010010111100010100100",
    737 => "10111111100101101100110000011010",
    738 => "10111111011011001010101110011111",
    739 => "00000000000000000000000000000000",
    740 => "00111111100000000000000000000000",
    741 => "00111110110001011100100001110101",
    742 => "00000000000000000000000000000000",
    743 => "00111101000100110000100101010001",
    744 => "10111110000000000000101101110001",
    745 => "00111111011010100001101110110101",
    746 => "00111111110010010000111111011000",
    747 => "00111111100000000000000000000000",
    748 => "00111111001110010110011111011000",
    749 => "00111111110010010000111111011000",
    750 => "00111111010000101110000101001011",
    751 => "00111111001100001001101001100111",
    752 => "00111101000000111010000000110001",
    753 => "10111101111011011001100001110000",
    754 => "00111111010110010100101111111101",
    755 => "10111111010000000001110100001010",
    756 => "10111111001011101001011011010110",
    757 => "00000000000000000000000000000000",
    758 => "00111111100000000000000000000000",
    759 => "00111111001110110100110000110011",
    760 => "00000000000000000000000000000000",
    761 => "00111101000001001000000110111001",
    762 => "10111101111011101011010010010010",
    763 => "00111111010110100101000011100110",
    764 => "00111111010000010000011111011110",
    765 => "00111111001011110100001001011011",
    766 => "00111111100000000000000000000000",
    767 => "00111111001110101010110000111000",
    768 => "00111101000001000111001001110101",
    769 => "10111101111011101010000101100100",
    770 => "00111111010110100011111101001100",
    771 => "10111111010000001111100000000101",
    772 => "10111111001011110011011011001101",
    773 => "00000000000000000000000000000000",
    774 => "00111111100000000000000000000000",
    775 => "00111111001110101011011100001000",
    776 => "00000000000000000000000000000000",
    777 => "00111101000001000111001101111001",
    778 => "10111101111011101010001010101011",
    779 => "00111111010110100100000001111000",
    780 => "00111111010000001111100100010101",
    781 => "00111111001011110011011110010011",
    782 => "00111111100000000000000000000000",
    783 => "00111111001110101011011001001101",
    784 => "00111101000001000111001101100010",
    785 => "10111101111011101010001010001110",
    786 => "00111111010110100100000001011101",
    787 => "10111111010000001111100011111010",
    788 => "10111111001011110011011101111111",
    789 => "00000000000000000000000000000000",
    790 => "00111111100000000000000000000000",
    791 => "00111111001110101011011001100000",
    792 => "00000000000000000000000000000000",
    793 => "00111101000001000111001101101010",
    794 => "10111101111011101010001010010111",
    795 => "00111111010110100100000001100110",
    796 => "00111111010000001111100100000101",
    797 => "00111111001011110011011110000111",
    798 => "00111111100000000000000000000000",
    799 => "00111111001110101011011001011001",
    800 => "00111101000001000111001101101000",
    801 => "10111101111011101010001010010101",
    802 => "00111111010110100100000001100101",
    803 => "10111111010000001111100100000001",
    804 => "10111111001011110011011110000100",
    805 => "00000000000000000000000000000000",
    806 => "00111111100000000000000000000000",
    807 => "00111111001110101011011001011100",
    808 => "00000000000000000000000000000000",
    809 => "00111101000001000111001101101000",
    810 => "10111101111011101010001010010101",
    811 => "00111111010110100100000001100101",
    812 => "00111111010000001111100100000011",
    813 => "00111111001011110011011110000110",
    814 => "00111111100000000000000000000000",
    815 => "00111111001110101011011001011010",
    816 => "00000000000000000000000000000000",
    817 => "00000000000000000000000000000000",
    818 => "00000000000000000000000000000000",
    819 => "00111101110000000010001000111101",
    820 => "10111110000100110001011000100111",
    821 => "00111111101010010111100010100100",
    822 => "00111110000001100000101011000010",
    823 => "00111110000001011010100011011000",
    824 => "00111111100000000000000000000000",
    825 => "00111111011111011100111101010011",
    826 => "00111101101111100111110101101111",
    827 => "10111110000101000110011110101011",
    828 => "00111111101010000010011010100001",
    829 => "00111111110010010000111111011000",
    830 => "00111111100000000000000000000000",
    831 => "00111111011010111001100001111101",
    832 => "00111111110010010000111111011000",
    833 => "00111110110011011100111111001000",
    834 => "00111110110010000101000001010010",
    835 => "00111101000101010011111110011000",
    836 => "10111110000000010100101010110010",
    837 => "00111111011011000101100000010001",
    838 => "00111101101110100000000101011000",
    839 => "00111101101110011011111111101000",
    840 => "00111111100000000000000000000000",
    841 => "00111111011111101111000111100100",
    842 => "00111101101110110000111101011000",
    843 => "10111110000101110000001101001011",
    844 => "00111111101001011010010110001001",
    845 => "00111111110010010000111111011000",
    846 => "00111111100000000000000000000000",
    847 => "00111111011010011100101111001100",
    848 => "00111111110010010000111111011000",
    849 => "00111110110101101101001110111000",
    850 => "00111110110100001001010000111111",
    851 => "00111101000110010001001010010111",
    852 => "10111110000000110110011001111010",
    853 => "00111111011100000001101010111101",
    854 => "00111101101111010000001101111011",
    855 => "00111101101111001011111011010001",
    856 => "00111111100000000000000000000000",
    857 => "00111111011111101110100100010110",
    858 => "00111101101110110010011000001000",
    859 => "10111110000101101111001010101011",
    860 => "00111111101001011011010100001110",
    861 => "00111111110010010000111111011000",
    862 => "00111111100000000000000000000000",
    863 => "00111111011010011101011100101011",
    864 => "00111111110010010000111111011000",
    865 => "00111110110101101001101111011100",
    866 => "00111110110100000110000100111010",
    867 => "00111101000110001111110001101110",
    868 => "10111110000000110101101001101110",
    869 => "00111111011100000000010101010010",
    870 => "00111101101111001111001001011001",
    871 => "00111101101111001010110111000001",
    872 => "00111111100000000000000000000000",
    873 => "00111111011111101110100101001000",
    874 => "00111101101110110010010110000011",
    875 => "10111110000101101111001100001100",
    876 => "00111111101001011011010010110110",
    877 => "00111111110010010000111111011000",
    878 => "00111111100000000000000000000000",
    879 => "00111111011010011101011011101011",
    880 => "00111111110010010000111111011000",
    881 => "00111110110101101001110100011000",
    882 => "00111110110100000110001001011010",
    883 => "00111101000110001111110011101011",
    884 => "10111110000000110101101010110010",
    885 => "00111111011100000000010111001100",
    886 => "00111101101111001111001010111011",
    887 => "00111101101111001010111000100011",
    888 => "00111111100000000000000000000000",
    889 => "00111111011111101110100101001000",
    890 => "00111101101110110010010110000111",
    891 => "10111110000101101111001100001001",
    892 => "00111111101001011011010010110111",
    893 => "00111111110010010000111111011000",
    894 => "00111111100000000000000000000000",
    895 => "00111111011010011101011011101011",
    896 => "00111111110010010000111111011000",
    897 => "00111110110101101001110100010100",
    898 => "00111110110100000110001001010111",
    899 => "00000000000000000000000000000000",
    900 => "00000000000000000000000000000000",
    901 => "00000000000000000000000000000000",
    902 => "00111111110011001100110011001110",
    903 => "00111111010011001100110011001110",
    904 => "00111101110000000010001000111101",
    905 => "10111110000100110001011000100111",
    906 => "00111111101010010111100010100100",
    907 => "10111110000001100000101010111010",
    908 => "10111110000001011010100011010000",
    909 => "00000000000000000000000000000000",
    910 => "00111111100000000000000000000000",
    911 => "00111111011111011100111101010011",
    912 => "00000000000000000000000000000000",
    913 => "00111101101111100111110101101111",
    914 => "10111110000101000110011110101011",
    915 => "00111111101010000010011010100001",
    916 => "00111111110010010000111111011000",
    917 => "00111111100000000000000000000000",
    918 => "00111111010010011111111110001100",
    919 => "00111111110010010000111111011000",
    920 => "00111111001010010110011000010000",
    921 => "00111111000111010100111010011000",
    922 => "00111101011010101101101101101110",
    923 => "10111110001000100001011010111111",
    924 => "00111111100100011001011000011101",
    925 => "10111101111001011101111000111000",
    926 => "10111101111001010110001010111110",
    927 => "00000000000000000000000000000000",
    928 => "00111111100000000000000000000000",
    929 => "00111111011111100110001110100001",
    930 => "00000000000000000000000000000000",
    931 => "00111101101111001111001010001011",
    932 => "10111110000101011001101000001011",
    933 => "00111111101001101111101111100011",
    934 => "00111111110010010000111111011000",
    935 => "00111111100000000000000000000000",
    936 => "00111111010010001111110111110100",
    937 => "00111111110010010000111111011000",
    938 => "00111111001010110000100001001100",
    939 => "00111111000111101001011111001000",
    940 => "00111101011010111001100000110000",
    941 => "10111110001000100011110110000111",
    942 => "00111111100100011011010100100100",
    943 => "10111101111001100000111111011101",
    944 => "10111101111001011001010000010010",
    945 => "00000000000000000000000000000000",
    946 => "00111111100000000000000000000000",
    947 => "00111111011111100110001011101110",
    948 => "00000000000000000000000000000000",
    949 => "00111101101111001111011000101100",
    950 => "10111110000101011001011101000110",
    951 => "00111111101001101111111010001110",
    952 => "00111111110010010000111111011000",
    953 => "00111111100000000000000000000000",
    954 => "00111111010010010000000001000011",
    955 => "00111111110010010000111111011000",
    956 => "00111111001010110000010010010000",
    957 => "00111111000111101001010011011010",
    958 => "00111101011010111001011010010111",
    959 => "10111110001000100011110100110100",
    960 => "00111111100100011011010011100010",
    961 => "10111101111001100000111101110011",
    962 => "10111101111001011001001110101001",
    963 => "00000000000000000000000000000000",
    964 => "00111111100000000000000000000000",
    965 => "00111111011111100110001011101111",
    966 => "00000000000000000000000000000000",
    967 => "00111101101111001111011000100100",
    968 => "10111110000101011001011101001100",
    969 => "00111111101001101111111010001001",
    970 => "00111111110010010000111111011000",
    971 => "00111111100000000000000000000000",
    972 => "00111111010010010000000000111110",
    973 => "00111111110010010000111111011000",
    974 => "00111111001010110000010010010111",
    975 => "00111111000111101001010011100000",
    976 => "00111101011010111001011010011011",
    977 => "10111110001000100011110100110101",
    978 => "00111111100100011011010011100010",
    979 => "10111101111001100000111101110011",
    980 => "10111101111001011001001110101001",
    981 => "00000000000000000000000000000000",
    982 => "00111111100000000000000000000000",
    983 => "00111111011111100110001011101111",
    984 => "00000000000000000000000000000000",
    985 => "00111101101111001111011000100100",
    986 => "10111110000101011001011101001100",
    987 => "00111111101001101111111010001001",
    988 => "00111111110010010000111111011000",
    989 => "00111111100000000000000000000000",
    990 => "00111111010010010000000000111110",
    991 => "00111111110010010000111111011000",
    992 => "00111111001010110000010010010111",
    993 => "00111111000111101001010011100000",
    994 => "00000000000000000000000000000000",
    995 => "00000000000000000000000000000000",
    996 => "00000000000000000000000000000000",
    997 => "00111101110000000010001000111101",
    998 => "10111110000100110001011000100111",
    999 => "00111111101010010111100010100100");

  constant b_lut : lut := (
    0 => "00111101011110011000100011001000",
    1 => "00110110001001100100110110101100",
    2 => "00111011111010000100011000001101",
    3 => "00110100000001001110000100001101",
    4 => "00111110000011000101110011110000",
    5 => "00110111111011001100100110010111",
    6 => "00111100110000111111101100011010",
    7 => "00110110000011011110010111010011",
    8 => "00111110111111111111111100000000",
    9 => "00111110101011110001110010001100",
    10 => "00111111011100001000111111010100",
    11 => "01000010101110111110111110100001",
    12 => "11000010100010001100111001001101",
    13 => "01000011001000101100001010111101",
    14 => "00111111010111110110010111111110",
    15 => "00111110011110011000110110000110",
    16 => "00111001001001100101011100101001",
    17 => "00111111010001000001101011100100",
    18 => "00111111010111110110010111111110",
    19 => "00111101011010000100110010101101",
    20 => "00110111100001001110100111100110",
    21 => "00111111010111110110010111111110",
    22 => "00111110011110011000110110000110",
    23 => "00111001001001100101011100101001",
    24 => "00111111010111110110010111111110",
    25 => "00111101011010000100110010101101",
    26 => "00110111100001001110100111100110",
    27 => "00111111000011100000000011010110",
    28 => "00111111100000000000000000000000",
    29 => "00111111011001100110011001100110",
    30 => "00111110000011101001010001101000",
    31 => "00111100100011110101001111000101",
    32 => "00111100011101011001100010011110",
    33 => "10111001110000111111111001110010",
    34 => "10101111000011011110101101111001",
    35 => "10111110000001011010100011011000",
    36 => "00111100000011000101111010001000",
    37 => "00110001111011001101000110101001",
    38 => "00111111011111011100111101010011",
    39 => "00111110000011101001010001101000",
    40 => "00111100100011110101001111000101",
    41 => "00111100011101011001100010011110",
    42 => "00111111100101011001101111100110",
    43 => "00111101101001010111011001101111",
    44 => "00110110110000011111000011111001",
    45 => "00111111100101011001101111100110",
    46 => "00111100001100010101110110011011",
    47 => "00110100101100100111010000101011",
    48 => "00111110000011101001010001101000",
    49 => "00111100100011110101001111000101",
    50 => "00111100011101011001100010011110",
    51 => "10111001000000101110110111000111",
    52 => "10101101001011111100010011100110",
    53 => "10111101101110011011111111101000",
    54 => "00111011100001110010010111110100",
    55 => "00110000010100110101110101001010",
    56 => "00111111011111101111000111100100",
    57 => "00111110000011101001010001101000",
    58 => "00111100100011110101001111000101",
    59 => "00111100011101011001100010011110",
    60 => "00111111100100110101101011101010",
    61 => "00111101101101000100011010100111",
    62 => "00110110111110101101010100101100",
    63 => "00111111100100110101101011101010",
    64 => "00111100010010011011010110100100",
    65 => "00110100111100001110100110000000",
    66 => "00111110000011101001010001101000",
    67 => "00111100100011110101001111000101",
    68 => "00111100011101011001100010011110",
    69 => "10111001000010010110001010000100",
    70 => "10101101010001001010100100100010",
    71 => "10111101101111001011111011010001",
    72 => "00111011100010111000111000100100",
    73 => "00110000011010001011100100001011",
    74 => "00111111011111101110100100010110",
    75 => "00111110000011101001010001101000",
    76 => "00111100100011110101001111000101",
    77 => "00111100011101011001100010011110",
    78 => "00111111100100110110100011100001",
    79 => "00111101101100111110100011110011",
    80 => "00110110111110010100111011010101",
    81 => "00111111100100110110100011100001",
    82 => "00111100010010010001100001110011",
    83 => "00110100111011110011010001010111",
    84 => "00111110000011101001010001101000",
    85 => "00111100100011110101001111000101",
    86 => "00111100011101011001100010011110",
    87 => "10111001000010010011110100101100",
    88 => "10101101010001000010110001111100",
    89 => "10111101101111001010110111000001",
    90 => "00111011100010110111010011011001",
    91 => "00110000011010000011101010010101",
    92 => "00111111011111101110100101001000",
    93 => "00111110000011101001010001101000",
    94 => "00111100100011110101001111000101",
    95 => "00111100011101011001100010011110",
    96 => "00111111100100110110100010010010",
    97 => "00111101101100111110101100000101",
    98 => "00110110111110010101011101110001",
    99 => "00111111100100110110100010010010",
    100 => "00111100010010010001101111101100",
    101 => "00110100111011110011110111111000",
    102 => "00111110000011101001010001101000",
    103 => "00111100100011110101001111000101",
    104 => "00111100011101011001100010011110",
    105 => "10111001000010010011111000000010",
    106 => "10101101010001000010111101000010",
    107 => "10111101101111001010111000100011",
    108 => "00111011100010110111010101101001",
    109 => "00110000011010000011110101101001",
    110 => "00111111011111101110100101001000",
    111 => "00111110000011101001010001101000",
    112 => "00111100100011110101001111000101",
    113 => "00111100011101011001100010011110",
    114 => "00111111100100110110100010010011",
    115 => "00111101101100111110101011111110",
    116 => "00110110111110010101011101010011",
    117 => "00111111100100110110100010010011",
    118 => "00111100010010010001101111100001",
    119 => "00110100111011110011110111011000",
    120 => "00111111000101100111110100111110",
    121 => "10111101011100101101101011101100",
    122 => "00111111010011101000101000101010",
    123 => "00111110000011101001010001101000",
    124 => "00111100100011110101001111000101",
    125 => "00111100011101011001100010011110",
    126 => "00111111100101101100110000011010",
    127 => "00111101100111011110100010000011",
    128 => "00110110101010001001001001100010",
    129 => "00111111100101101100110000011010",
    130 => "00111100001001010101101111001101",
    131 => "00110100100101111000011100101010",
    132 => "00111110000011101001010001101000",
    133 => "00111100100011110101001111000101",
    134 => "00111100011101011001100010011110",
    135 => "00111111010011110100000110101101",
    136 => "00111110100101000101010100111110",
    137 => "00111001100010111011101001100000",
    138 => "00111111010011110100000110101101",
    139 => "00111101100101101000110001100011",
    140 => "00110111111100110111011100111100",
    141 => "00111110000011101001010001101000",
    142 => "00111100100011110101001111000101",
    143 => "00111100011101011001100010011110",
    144 => "00111101100100000100000100010110",
    145 => "00110111110111000101111111000001",
    146 => "00111110100100000010101101010101",
    147 => "00111001100000000100100111101100",
    148 => "00111110000011101001010001101000",
    149 => "00111100100011110101001111000101",
    150 => "00111100011101011001100010011110",
    151 => "00111101100100100101010011111100",
    152 => "00110111111000111101100111111000",
    153 => "00111110100100011000110011100000",
    154 => "00111001100001000000001011001010",
    155 => "00111110000011101001010001101000",
    156 => "00111100100011110101001111000101",
    157 => "00111100011101011001100010011110",
    158 => "00111101100100100011000011110000",
    159 => "00110111111000110101011100011001",
    160 => "00111110100100010111010011111001",
    161 => "00111001100000111100000111001001",
    162 => "00111110000011101001010001101000",
    163 => "00111100100011110101001111000101",
    164 => "00111100011101011001100010011110",
    165 => "00111101100100100011001101010110",
    166 => "00110111111000110101111111001110",
    167 => "00111110100100010111011010010000",
    168 => "00111001100000111100011000011011",
    169 => "00111110000011101001010001101000",
    170 => "00111100100011110101001111000101",
    171 => "00111100011101011001100010011110",
    172 => "00111101100100100011001100101011",
    173 => "00110111111000110101111100110000",
    174 => "00111110100100010111011001110011",
    175 => "00111001100000111100010111001101",
    176 => "00111110000011101001010001101000",
    177 => "00111100100011110101001111000101",
    178 => "00111100011101011001100010011110",
    179 => "00111101100100100011001100110010",
    180 => "00110111111000110101111101001000",
    181 => "00111110100100010111011001110111",
    182 => "00111001100000111100010111011001",
    183 => "00111110000011101001010001101000",
    184 => "00111100100011110101001111000101",
    185 => "00111100011101011001100010011110",
    186 => "00111101100100100011001100101011",
    187 => "00110111111000110101111100110000",
    188 => "00111110100100010111011001110011",
    189 => "00111001100000111100010111001101",
    190 => "00111110000011101001010001101000",
    191 => "00111100100011110101001111000101",
    192 => "00111100011101011001100010011110",
    193 => "00111101100100100011001100110010",
    194 => "00110111111000110101111101001000",
    195 => "00111110100100010111011001110111",
    196 => "00111001100000111100010111011001",
    197 => "00111111000010111110011110000001",
    198 => "00111111000010111110011101111111",
    199 => "00111111001000100111001011100000",
    200 => "00111111011001100110011001100110",
    201 => "00111110000011101001010001101000",
    202 => "00111100100011110101001111000101",
    203 => "00111100011101011001100010011110",
    204 => "10111100001001010101111010101101",
    205 => "10110100100101111000110101001101",
    206 => "10111110110000111110111101010110",
    207 => "00111101100111011110101001010111",
    208 => "00110110101010001001100000111101",
    209 => "00111111011011001000001101010001",
    210 => "00111110000011101001010001101000",
    211 => "00111100100011110101001111000101",
    212 => "00111100011101011001100010011110",
    213 => "00111111100011100111101001000101",
    214 => "00111101110101101000000111100001",
    215 => "00110111010100110100100010111101",
    216 => "00111111100011100111101001000101",
    217 => "00111100100000101110011101101010",
    218 => "00110101010111010101101101101100",
    219 => "00111110000011101001010001101000",
    220 => "00111100100011110101001111000101",
    221 => "00111100011101011001100010011110",
    222 => "10111011011110010001010001111100",
    223 => "10110010111110000100011010011000",
    224 => "10111110100011110100000010111101",
    225 => "00111101001001001011000011011101",
    226 => "00110101001111110011110101111010",
    227 => "00111111011101011100011010001110",
    228 => "00111110000011101001010001101000",
    229 => "00111100100011110101001111000101",
    230 => "00111100011101011001100010011110",
    231 => "00111111100010001100011000101111",
    232 => "00111110000000010010011101001111",
    233 => "00110111101110000111011110100000",
    234 => "00111111100010001100011000101111",
    235 => "00111100101011001111101010110010",
    236 => "00110101110101000001001110100101",
    237 => "00111110000011101001010001101000",
    238 => "00111100100011110101001111000101",
    239 => "00111100011101011001100010011110",
    240 => "10111011011101000011111111100111",
    241 => "10110010111011010010111110101100",
    242 => "10111110100011100101100001111110",
    243 => "00111101001000101000111000000010",
    244 => "00110101001101111110010100001001",
    245 => "00111111011101011110100001001000",
    246 => "00111110000011101001010001101000",
    247 => "00111100100011110101001111000101",
    248 => "00111100011101011001100010011110",
    249 => "00111111100010001011110010011000",
    250 => "00111110000000010100110111011010",
    251 => "00110111101110010001110011111000",
    252 => "00111111100010001011110010011000",
    253 => "00111100101011010100100000100101",
    254 => "00110101110101001111000101111011",
    255 => "00111110000011101001010001101000",
    256 => "00111100100011110101001111000101",
    257 => "00111100011101011001100010011110",
    258 => "10111011011101000000010110111110",
    259 => "10110010111011001010101111110111",
    260 => "10111110100011100100110101111111",
    261 => "00111101001000100111010000110011",
    262 => "00110101001101111000110110000001",
    263 => "00111111011101011110100111100000",
    264 => "00111110000011101001010001101000",
    265 => "00111100100011110101001111000101",
    266 => "00111100011101011001100010011110",
    267 => "00111111100010001011110000100101",
    268 => "00111110000000010100111110101000",
    269 => "00110111101110010010010010111010",
    270 => "00111111100010001011110000100101",
    271 => "00111100101011010100101111000111",
    272 => "00110101110101001111101111100100",
    273 => "00111110000011101001010001101000",
    274 => "00111100100011110101001111000101",
    275 => "00111100011101011001100010011110",
    276 => "10111011011101000000001100001101",
    277 => "10110010111011001010010111100001",
    278 => "10111110100011100100110011111011",
    279 => "00111101001000100111001100000001",
    280 => "00110101001101111000100101110010",
    281 => "00111111011101011110100111110010",
    282 => "00111110000011101001010001101000",
    283 => "00111100100011110101001111000101",
    284 => "00111100011101011001100010011110",
    285 => "00111111100010001011110000100000",
    286 => "00111110000000010100111110111100",
    287 => "00110111101110010010010100001111",
    288 => "00111111100010001011110000100000",
    289 => "00111100101011010100101111110000",
    290 => "00110101110101001111110001011010",
    291 => "00111111000100010000100001100001",
    292 => "10111110001101111111110000110011",
    293 => "00111111010011011110000011010100",
    294 => "00111110000011101001010001101000",
    295 => "00111100100011110101001111000101",
    296 => "00111100011101011001100010011110",
    297 => "00111111011010101001001011010101",
    298 => "00111110010110110101001000101000",
    299 => "00111000111000011101010001010111",
    300 => "00111111011010101001001011010101",
    301 => "00111101001111110110010001110100",
    302 => "00110111001010010010101001001101",
    303 => "00111110000011101001010001101000",
    304 => "00111100100011110101001111000101",
    305 => "00111100011101011001100010011110",
    306 => "00111111100000010010100101000010",
    307 => "00111110001000011000110110111000",
    308 => "00111000001101001000010010010110",
    309 => "00111111100000010010100101000010",
    310 => "00111100111100011111111100101010",
    311 => "00110110011010000001110011100010",
    312 => "00111110000011101001010001101000",
    313 => "00111100100011110101001111000101",
    314 => "00111100011101011001100010011110",
    315 => "00111101000101001100111100010110",
    316 => "00110110101111000001000111000000",
    317 => "00111110001110010111001000001101",
    318 => "00111000100010001000010010010001",
    319 => "00111110000011101001010001101000",
    320 => "00111100100011110101001111000101",
    321 => "00111100011101011001100010011110",
    322 => "00111111011001110111110111000110",
    323 => "00111110011000110111011011100100",
    324 => "00111000111110111110111000111001",
    325 => "00111111011001110111110111000110",
    326 => "00111101010010100010011010000100",
    327 => "00110111010000000011000001010011",
    328 => "00111110000011101001010001101000",
    329 => "00111100100011110101001111000101",
    330 => "00111100011101011001100010011110",
    331 => "00111101000001101110100010001001",
    332 => "00110110100101011001101001101010",
    333 => "00111110001011011011010110001110",
    334 => "00111000011000000110100010000110",
    335 => "00111110000011101001010001101000",
    336 => "00111100100011110101001111000101",
    337 => "00111100011101011001100010011110",
    338 => "00111111011001110000111011110101",
    339 => "00111110011001001001111010110111",
    340 => "00111000111111111100101000101011",
    341 => "00111111011001110000111011110101",
    342 => "00111101010010111011000101100001",
    343 => "00110111010000111010000010111001",
    344 => "00111110000011101001010001101000",
    345 => "00111100100011110101001111000101",
    346 => "00111100011101011001100010011110",
    347 => "00111101000001101101111111101010",
    348 => "00110110100101011000010000011110",
    349 => "00111110001011011010111000101000",
    350 => "00111000011000000100101111011010",
    351 => "00111110000011101001010001101000",
    352 => "00111100100011110101001111000101",
    353 => "00111100011101011001100010011110",
    354 => "00111111011001110000111010111010",
    355 => "00111110011001001001111101010101",
    356 => "00111000111111111100110000111010",
    357 => "00111111011001110000111010111010",
    358 => "00111101010010111011001000110010",
    359 => "00110111010000111010001010010001",
    360 => "00111110000011101001010001101000",
    361 => "00111100100011110101001111000101",
    362 => "00111100011101011001100010011110",
    363 => "00111101000001101101111111100010",
    364 => "00110110100101011000010000001000",
    365 => "00111110001011011010111000100001",
    366 => "00111000011000000100101111000000",
    367 => "00111110000011101001010001101000",
    368 => "00111100100011110101001111000101",
    369 => "00111100011101011001100010011110",
    370 => "00111111011001110000111010110110",
    371 => "00111110011001001001111101100000",
    372 => "00111000111111111100110001011110",
    373 => "00111111011001110000111010110110",
    374 => "00111101010010111011001001000010",
    375 => "00110111010000111010001010110000",
    376 => "00111111000110001010111000000001",
    377 => "00111110110101011111110011001000",
    378 => "00111111001011110110111100111100",
    379 => "00111111011001100110011001100110",
    380 => "00111110000011101001010001101000",
    381 => "00111100100011110101001111000101",
    382 => "00111100011101011001100010011110",
    383 => "10111101001111110110011001110101",
    384 => "10110111001010010010111001110010",
    385 => "10111111000110111101011111111000",
    386 => "00111110010110110101001110110001",
    387 => "00111000111000011101100100010111",
    388 => "00111111010010110001100100010011",
    389 => "00111110000011101001010001101000",
    390 => "00111100100011110101001111000101",
    391 => "00111100011101011001100010011110",
    392 => "00111111100001111111011110101111",
    393 => "00111110000001000110101000111010",
    394 => "00110111110001101100110000111010",
    395 => "00111111100001111111011110101111",
    396 => "00111100101100111001001010010111",
    397 => "00110101111001110110101101110110",
    398 => "00111110000011101001010001101000",
    399 => "00111100100011110101001111000101",
    400 => "00111100011101011001100010011110",
    401 => "10111100100010100000011100111111",
    402 => "10110101011110100111111001000100",
    403 => "10111110111001011111101011010011",
    404 => "00111101110111100011100010101001",
    405 => "00110111011010101110100001101100",
    406 => "00111111011001001011100010010111",
    407 => "00111110000011101001010001101000",
    408 => "00111100100011110101001111000101",
    409 => "00111100011101011001100010011110",
    410 => "00111111100000100010011100000000",
    411 => "00111110000111010010000101010001",
    412 => "00111000001001100001011110010010",
    413 => "00111111100000100010011100000000",
    414 => "00111100111010000010000001000010",
    415 => "00110110010100101001111010101010",
    416 => "00111110000011101001010001101000",
    417 => "00111100100011110101001111000101",
    418 => "00111100011101011001100010011110",
    419 => "10111100010111011010101010100010",
    420 => "10110101000101100001111001010000",
    421 => "10111110110101101101001111110011",
    422 => "00111101101111111111101010011111",
    423 => "00110111000101110111011000010110",
    424 => "00111111011010000110000000001110",
    425 => "00111110000011101001010001101000",
    426 => "00111100100011110101001111000101",
    427 => "00111100011101011001100010011110",
    428 => "00111111100000011001001101111011",
    429 => "00111110000111111011000111000001",
    430 => "00111000001011100101101101011111",
    431 => "00111111100000011001001101111011",
    432 => "00111100111011011101010011001100",
    433 => "00110110010111101110010110101010",
    434 => "00111110000011101001010001101000",
    435 => "00111100100011110101001111000101",
    436 => "00111100011101011001100010011110",
    437 => "10111100010110101100100101101011",
    438 => "10110101000100011001101101110011",
    439 => "10111110110101011111001111001100",
    440 => "00111101101111100101000000001011",
    441 => "00110111000100111000110100101110",
    442 => "00111111011010001001001110111100",
    443 => "00111110000011101001010001101000",
    444 => "00111100100011110101001111000101",
    445 => "00111100011101011001100010011110",
    446 => "00111111100000011000101111110101",
    447 => "00111110000111111101001101100000",
    448 => "00111000001011101100100110010101",
    449 => "00111111100000011000101111110101",
    450 => "00111100111011100001111111101011",
    451 => "00110110010111111000101000010000",
    452 => "00111110000011101001010001101000",
    453 => "00111100100011110101001111000101",
    454 => "00111100011101011001100010011110",
    455 => "10111100010110101010011000011110",
    456 => "10110101000100010110010010100110",
    457 => "10111110110101011110100100000010",
    458 => "00111101101111100011101110010001",
    459 => "00110111000100110101110110010011",
    460 => "00111111011010001001011000110111",
    461 => "00111110000011101001010001101000",
    462 => "00111100100011110101001111000101",
    463 => "00111100011101011001100010011110",
    464 => "00111111100000011000101110011010",
    465 => "00111110000111111101010011110111",
    466 => "00111000001011101100111011001100",
    467 => "00111111100000011000101110011010",
    468 => "00111100111011100010001101111001",
    469 => "00110110010111111001000111011000",
    470 => "00111111000110110001111110000110",
    471 => "10111110100110001101110011011001",
    472 => "00111111001111001100001100010000",
    473 => "00111110000011101001010001101000",
    474 => "00111100100011110101001111000101",
    475 => "00111100011101011001100010011110",
    476 => "00111101001111110110011010000000",
    477 => "00110111001010010010111010000101",
    478 => "00111110010110110101001110111000",
    479 => "00111000111000011101100100101101",
    480 => "00111110000011101001010001101000",
    481 => "00111100100011110101001111000101",
    482 => "00111100011101011001100010011110",
    483 => "00111111100001111111011110101111",
    484 => "00111110000001000110101000111010",
    485 => "00110111110001101100110000111010",
    486 => "00111111100001111111011110101111",
    487 => "00111100101100111001001010010111",
    488 => "00110101111001110110101101110110",
    489 => "00111110000011101001010001101000",
    490 => "00111100100011110101001111000101",
    491 => "00111100011101011001100010011110",
    492 => "00111100100010100000011101000100",
    493 => "00110101011110100111111001011010",
    494 => "00111101110111100011100010101110",
    495 => "00110111011010101110100010000000",
    496 => "00111110000011101001010001101000",
    497 => "00111100100011110101001111000101",
    498 => "00111100011101011001100010011110",
    499 => "00111111100000100010011011111111",
    500 => "00111110000111010010000101010101",
    501 => "00111000001001100001011110011111",
    502 => "00111111100000100010011011111111",
    503 => "00111100111010000010000001001011",
    504 => "00110110010100101001111010111111",
    505 => "00111110000011101001010001101000",
    506 => "00111100100011110101001111000101",
    507 => "00111100011101011001100010011110",
    508 => "00111100010111011010101010101011",
    509 => "00110101000101100001111001011111",
    510 => "00111101101111111111101010100101",
    511 => "00110111000101110111011000100011",
    512 => "00111110000011101001010001101000",
    513 => "00111100100011110101001111000101",
    514 => "00111100011101011001100010011110",
    515 => "00111111100000011001001101111100",
    516 => "00111110000111111011000110111101",
    517 => "00111000001011100101101101010000",
    518 => "00111111100000011001001101111100",
    519 => "00111100111011011101010011000010",
    520 => "00110110010111101110010110010010",
    521 => "00111110000011101001010001101000",
    522 => "00111100100011110101001111000101",
    523 => "00111100011101011001100010011110",
    524 => "00111100010110101100100101101111",
    525 => "00110101000100011001101101111000",
    526 => "00111101101111100101000000001101",
    527 => "00110111000100111000110100110011",
    528 => "00111110000011101001010001101000",
    529 => "00111100100011110101001111000101",
    530 => "00111100011101011001100010011110",
    531 => "00111111100000011000101111110100",
    532 => "00111110000111111101001101100100",
    533 => "00111000001011101100100110100010",
    534 => "00111111100000011000101111110100",
    535 => "00111100111011100001111111110101",
    536 => "00110110010111111000101000100110",
    537 => "00111110000011101001010001101000",
    538 => "00111100100011110101001111000101",
    539 => "00111100011101011001100010011110",
    540 => "00111100010110101010011000100111",
    541 => "00110101000100010110010010110100",
    542 => "00111101101111100011101110010110",
    543 => "00110111000100110101110110011101",
    544 => "00111110000011101001010001101000",
    545 => "00111100100011110101001111000101",
    546 => "00111100011101011001100010011110",
    547 => "00111111100000011000101110011010",
    548 => "00111110000111111101010011110111",
    549 => "00111000001011101100111011001100",
    550 => "00111111100000011000101110011010",
    551 => "00111100111011100010001101111001",
    552 => "00110110010111111001000111011000",
    553 => "00111111000110110001111110001000",
    554 => "00111110100110001101110011011100",
    555 => "00111111001111001100001100010000",
    556 => "00111111011001100110011001100110",
    557 => "00111110000011101001010001101000",
    558 => "00111100100011110101001111000101",
    559 => "00111100011101011001100010011110",
    560 => "10111110000000110100110011110011",
    561 => "10111000110111101110110011011100",
    562 => "10111111010010110001100101100000",
    563 => "00111110110101101111000010111111",
    564 => "00111010010101001001000100000010",
    565 => "00111111000110111101011101010110",
    566 => "00111110000011101001010001101000",
    567 => "00111100100011110101001111000101",
    568 => "00111100011101011001100010011110",
    569 => "00111111100000010010100100111110",
    570 => "00111110001000011000110111001010",
    571 => "00111000001101001000010011010010",
    572 => "00111111100000010010100100111110",
    573 => "00111100111100011111111101010001",
    574 => "00110110011010000001110100111100",
    575 => "00111110000011101001010001101000",
    576 => "00111100100011110101001111000101",
    577 => "00111100011101011001100010011110",
    578 => "10111101000101001100111100000101",
    579 => "10110110101111000001000110001101",
    580 => "10111111000100001110111101000010",
    581 => "00111110001110010111000111111110",
    582 => "00111000100010001000010001110000",
    583 => "00111111010100110000010101110000",
    584 => "00111110000011101001010001101000",
    585 => "00111100100011110101001111000101",
    586 => "00111100011101011001100010011110",
    587 => "00111111011001110111110111000100",
    588 => "00111110011000110111011011101001",
    589 => "00111000111110111110111001001011",
    590 => "00111111011001110111110111000100",
    591 => "00111101010010100010011010001100",
    592 => "00110111010000000011000001100100",
    593 => "00111110000011101001010001101000",
    594 => "00111100100011110101001111000101",
    595 => "00111100011101011001100010011110",
    596 => "10111101000001101110100010000011",
    597 => "10110110100101011001101001011011",
    598 => "10111111000011001101001011001001",
    599 => "00111110001011011011010110001001",
    600 => "00111000011000000110100001110100",
    601 => "00111111010101011100100101101001",
    602 => "00111110000011101001010001101000",
    603 => "00111100100011110101001111000101",
    604 => "00111100011101011001100010011110",
    605 => "00111111011001110000111011111001",
    606 => "00111110011001001001111010101101",
    607 => "00111000111111111100101000000110",
    608 => "00111111011001110000111011111001",
    609 => "00111101010010111011000101010010",
    610 => "00110111010000111010000010011010",
    611 => "00111110000011101001010001101000",
    612 => "00111100100011110101001111000101",
    613 => "00111100011101011001100010011110",
    614 => "10111101000001101101111111100101",
    615 => "10110110100101011000010000001111",
    616 => "10111111000011001101000000100011",
    617 => "00111110001011011010111000100011",
    618 => "00111000011000000100101111001000",
    619 => "00111111010101011100101100101000",
    620 => "00111110000011101001010001101000",
    621 => "00111100100011110101001111000101",
    622 => "00111100011101011001100010011110",
    623 => "00111111011001110000111010110110",
    624 => "00111110011001001001111101100000",
    625 => "00111000111111111100110001011110",
    626 => "00111111011001110000111010110110",
    627 => "00111101010010111011001001000010",
    628 => "00110111010000111010001010110000",
    629 => "00111110000011101001010001101000",
    630 => "00111100100011110101001111000101",
    631 => "00111100011101011001100010011110",
    632 => "10111101000001101101111111100101",
    633 => "10110110100101011000010000001111",
    634 => "10111111000011001101000000100011",
    635 => "00111110001011011010111000100011",
    636 => "00111000011000000100101111001000",
    637 => "00111111010101011100101100101000",
    638 => "00111110000011101001010001101000",
    639 => "00111100100011110101001111000101",
    640 => "00111100011101011001100010011110",
    641 => "00111111011001110000111010110110",
    642 => "00111110011001001001111101100000",
    643 => "00111000111111111100110001011110",
    644 => "00111111011001110000111010110110",
    645 => "00111101010010111011001001000010",
    646 => "00110111010000111010001010110000",
    647 => "00111111000110001010111000000001",
    648 => "10111110110101011111110011000110",
    649 => "00111111001011110110111100111110",
    650 => "00111110000011101001010001101000",
    651 => "00111100100011110101001111000101",
    652 => "00111100011101011001100010011110",
    653 => "00111100001001010101111010110010",
    654 => "00110100100101111000110101011000",
    655 => "00111101100111011110101001011010",
    656 => "00110110101010001001100001000110",
    657 => "00111110000011101001010001101000",
    658 => "00111100100011110101001111000101",
    659 => "00111100011101011001100010011110",
    660 => "00111111100011100111101001000101",
    661 => "00111101110101101000000111100001",
    662 => "00110111010100110100100010111101",
    663 => "00111111100011100111101001000101",
    664 => "00111100100000101110011101101010",
    665 => "00110101010111010101101101101100",
    666 => "00111110000011101001010001101000",
    667 => "00111100100011110101001111000101",
    668 => "00111100011101011001100010011110",
    669 => "00111011011110010001010010000100",
    670 => "00110010111110000100011010101110",
    671 => "00111101001001001011000011100010",
    672 => "00110101001111110011110110001001",
    673 => "00111110000011101001010001101000",
    674 => "00111100100011110101001111000101",
    675 => "00111100011101011001100010011110",
    676 => "00111111100010001100011000101111",
    677 => "00111110000000010010011101001111",
    678 => "00110111101110000111011110100000",
    679 => "00111111100010001100011000101111",
    680 => "00111100101011001111101010110010",
    681 => "00110101110101000001001110100101",
    682 => "00111110000011101001010001101000",
    683 => "00111100100011110101001111000101",
    684 => "00111100011101011001100010011110",
    685 => "00111011011101000011111111110010",
    686 => "00110010111011010010111111000010",
    687 => "00111101001000101000111000000110",
    688 => "00110101001101111110010100011000",
    689 => "00111110000011101001010001101000",
    690 => "00111100100011110101001111000101",
    691 => "00111100011101011001100010011110",
    692 => "00111111100010001011110010011000",
    693 => "00111110000000010100110111011010",
    694 => "00110111101110010001110011111000",
    695 => "00111111100010001011110010011000",
    696 => "00111100101011010100100000100101",
    697 => "00110101110101001111000101111011",
    698 => "00111110000011101001010001101000",
    699 => "00111100100011110101001111000101",
    700 => "00111100011101011001100010011110",
    701 => "00111011011101000000010111001010",
    702 => "00110010111011001010110000010001",
    703 => "00111101001000100111010000110111",
    704 => "00110101001101111000110110001111",
    705 => "00111110000011101001010001101000",
    706 => "00111100100011110101001111000101",
    707 => "00111100011101011001100010011110",
    708 => "00111111100010001011110000100101",
    709 => "00111110000000010100111110101000",
    710 => "00110111101110010010010010111010",
    711 => "00111111100010001011110000100101",
    712 => "00111100101011010100101111000111",
    713 => "00110101110101001111101111100100",
    714 => "00111110000011101001010001101000",
    715 => "00111100100011110101001111000101",
    716 => "00111100011101011001100010011110",
    717 => "00111011011101000000001100010111",
    718 => "00110010111011001010010111110101",
    719 => "00111101001000100111001100000101",
    720 => "00110101001101111000100110000001",
    721 => "00111110000011101001010001101000",
    722 => "00111100100011110101001111000101",
    723 => "00111100011101011001100010011110",
    724 => "00111111100010001011110000011111",
    725 => "00111110000000010100111111000000",
    726 => "00110111101110010010010100100010",
    727 => "00111111100010001011110000011111",
    728 => "00111100101011010100101111111000",
    729 => "00110101110101001111110001110001",
    730 => "00111111000100010000100001100010",
    731 => "00111110001101111111110000110110",
    732 => "00111111010011011110000011010100",
    733 => "00111111011001100110011001100110",
    734 => "00111110000011101001010001101000",
    735 => "00111100100011110101001111000101",
    736 => "00111100011101011001100010011110",
    737 => "10111110100010111000011111100011",
    738 => "10111010001000011101011010001010",
    739 => "10111111011011001000001100101001",
    740 => "00111111001100011010011110100100",
    741 => "00111011011100000000110011001000",
    742 => "00111110110000111110100001011100",
    743 => "00111110000011101001010001101000",
    744 => "00111100100011110101001111000101",
    745 => "00111100011101011001100010011110",
    746 => "00111111010011110011111001100101",
    747 => "00111110100101000101101000111100",
    748 => "00111001100010111100100001111111",
    749 => "00111111010011110011111001100101",
    750 => "00111101100101101001001111111110",
    751 => "00110111111100111001001111110011",
    752 => "00111110000011101001010001101000",
    753 => "00111100100011110101001111000101",
    754 => "00111100011101011001100010011110",
    755 => "10111101100100000100000101110011",
    756 => "10110111110111000110000100001001",
    757 => "10111111001011101001010100011101",
    758 => "00111110100100000010101110010011",
    759 => "00111001100000000100101010010000",
    760 => "00111111001110110011110000101010",
    761 => "00111110000011101001010001101000",
    762 => "00111100100011110101001111000101",
    763 => "00111100011101011001100010011110",
    764 => "00111101100100100101010011110111",
    765 => "00110111111000111101100111101001",
    766 => "00111110100100011000110011011101",
    767 => "00111001100001000000001011000011",
    768 => "00111110000011101001010001101000",
    769 => "00111100100011110101001111000101",
    770 => "00111100011101011001100010011110",
    771 => "10111101100100100011000011110000",
    772 => "10110111111000110101011100011001",
    773 => "10111111001011110011010100000110",
    774 => "00111110100100010111010011111001",
    775 => "00111001100000111100000111001001",
    776 => "00111111001110101010011010010000",
    777 => "00111110000011101001010001101000",
    778 => "00111100100011110101001111000101",
    779 => "00111100011101011001100010011110",
    780 => "00111101100100100011001101011011",
    781 => "00110111111000110101111111011011",
    782 => "00111110100100010111011010010011",
    783 => "00111001100000111100011000100100",
    784 => "00111110000011101001010001101000",
    785 => "00111100100011110101001111000101",
    786 => "00111100011101011001100010011110",
    787 => "10111101100100100011001100011110",
    788 => "10110111111000110101111011111101",
    789 => "10111111001011110011010110111000",
    790 => "00111110100100010111011001101010",
    791 => "00111001100000111100010110110100",
    792 => "00111111001110101010010111100111",
    793 => "00111110000011101001010001101000",
    794 => "00111100100011110101001111000101",
    795 => "00111100011101011001100010011110",
    796 => "00111101100100100011001100110110",
    797 => "00110111111000110101111101011000",
    798 => "00111110100100010111011001111010",
    799 => "00111001100000111100010111100001",
    800 => "00111110000011101001010001101000",
    801 => "00111100100011110101001111000101",
    802 => "00111100011101011001100010011110",
    803 => "10111101100100100011001100101101",
    804 => "10110111111000110101111100110111",
    805 => "10111111001011110011010110111101",
    806 => "00111110100100010111011001110100",
    807 => "00111001100000111100010111010001",
    808 => "00111111001110101010010111100011",
    809 => "00111110000011101001010001101000",
    810 => "00111100100011110101001111000101",
    811 => "00111100011101011001100010011110",
    812 => "00111101100100100011001100110010",
    813 => "00110111111000110101111101001000",
    814 => "00111110100100010111011001110111",
    815 => "00111001100000111100010111011001",
    816 => "00111111000010111110011110000001",
    817 => "10111111000010111110011101111110",
    818 => "00111111001000100111001011100000",
    819 => "00111110000011101001010001101000",
    820 => "00111100100011110101001111000101",
    821 => "00111100011101011001100010011110",
    822 => "00111001110000111111111001110010",
    823 => "00101111000011011110101101111001",
    824 => "00111100000011000101111010001000",
    825 => "00110001111011001101000110101001",
    826 => "00111110000011101001010001101000",
    827 => "00111100100011110101001111000101",
    828 => "00111100011101011001100010011110",
    829 => "00111111100101011001101111100110",
    830 => "00111101101001010111011001101111",
    831 => "00110110110000011111000011111001",
    832 => "00111111100101011001101111100110",
    833 => "00111100001100010101110110011011",
    834 => "00110100101100100111010000101011",
    835 => "00111110000011101001010001101000",
    836 => "00111100100011110101001111000101",
    837 => "00111100011101011001100010011110",
    838 => "00111001000000101110110111000111",
    839 => "00101101001011111100010011100110",
    840 => "00111011100001110010010111110100",
    841 => "00110000010100110101110101001010",
    842 => "00111110000011101001010001101000",
    843 => "00111100100011110101001111000101",
    844 => "00111100011101011001100010011110",
    845 => "00111111100100110101101011101010",
    846 => "00111101101101000100011010100111",
    847 => "00110110111110101101010100101100",
    848 => "00111111100100110101101011101010",
    849 => "00111100010010011011010110100100",
    850 => "00110100111100001110100110000000",
    851 => "00111110000011101001010001101000",
    852 => "00111100100011110101001111000101",
    853 => "00111100011101011001100010011110",
    854 => "00111001000010010110001010000100",
    855 => "00101101010001001010100100100010",
    856 => "00111011100010111000111000100100",
    857 => "00110000011010001011100100001011",
    858 => "00111110000011101001010001101000",
    859 => "00111100100011110101001111000101",
    860 => "00111100011101011001100010011110",
    861 => "00111111100100110110100011100001",
    862 => "00111101101100111110100011110011",
    863 => "00110110111110010100111011010101",
    864 => "00111111100100110110100011100001",
    865 => "00111100010010010001100001110011",
    866 => "00110100111011110011010001010111",
    867 => "00111110000011101001010001101000",
    868 => "00111100100011110101001111000101",
    869 => "00111100011101011001100010011110",
    870 => "00111001000010010011110100101100",
    871 => "00101101010001000010110001111100",
    872 => "00111011100010110111010011011001",
    873 => "00110000011010000011101010010101",
    874 => "00111110000011101001010001101000",
    875 => "00111100100011110101001111000101",
    876 => "00111100011101011001100010011110",
    877 => "00111111100100110110100010010010",
    878 => "00111101101100111110101100000101",
    879 => "00110110111110010101011101110001",
    880 => "00111111100100110110100010010010",
    881 => "00111100010010010001101111101100",
    882 => "00110100111011110011110111111000",
    883 => "00111110000011101001010001101000",
    884 => "00111100100011110101001111000101",
    885 => "00111100011101011001100010011110",
    886 => "00111001000010010011111000000010",
    887 => "00101101010001000010111101000010",
    888 => "00111011100010110111010101101001",
    889 => "00110000011010000011110101101001",
    890 => "00111110000011101001010001101000",
    891 => "00111100100011110101001111000101",
    892 => "00111100011101011001100010011110",
    893 => "00111111100100110110100010010011",
    894 => "00111101101100111110101011111110",
    895 => "00110110111110010101011101010011",
    896 => "00111111100100110110100010010011",
    897 => "00111100010010010001101111100001",
    898 => "00110100111011110011110111011000",
    899 => "00111111000101100111110100111110",
    900 => "00111101011100101101101011101100",
    901 => "00111111010011101000101000101010",
    902 => "00111111011001100110011001100110",
    903 => "00111111011001100110011001100110",
    904 => "00111110000011101001010001101000",
    905 => "00111100100011110101001111000101",
    906 => "00111100011101011001100010011110",
    907 => "10111001110000111111111001001111",
    908 => "10101111000011011110101100111101",
    909 => "10111110000001011010100011010000",
    910 => "00111100000011000101111001110111",
    911 => "00110001111011001101000101010101",
    912 => "00111111011111011100111101010011",
    913 => "00111110000011101001010001101000",
    914 => "00111100100011110101001111000101",
    915 => "00111100011101011001100010011110",
    916 => "00111111011010001011100110100000",
    917 => "00111110011000000010111111010101",
    918 => "00111000111100010011001001000110",
    919 => "00111111011010001011100110100000",
    920 => "00111101010001011100110000001001",
    921 => "00110111001101101010101101101110",
    922 => "00111110000011101001010001101000",
    923 => "00111100100011110101001111000101",
    924 => "00111100011101011001100010011110",
    925 => "10111001011101110001110011101001",
    926 => "10101110010000010111000111001001",
    927 => "10111101111001010110001010111110",
    928 => "00111011110011100110011101010010",
    929 => "00110001001111000011101101000001",
    930 => "00111111011111100110001110100001",
    931 => "00111110000011101001010001101000",
    932 => "00111100100011110101001111000101",
    933 => "00111100011101011001100010011110",
    934 => "00111111011001110001011101100100",
    935 => "00111110011001001000100000101101",
    936 => "00111000111111110111111010001001",
    937 => "00111111011001110001011101100100",
    938 => "00111101010010111001001101000010",
    939 => "00110111010000110101110101000001",
    940 => "00111110000011101001010001101000",
    941 => "00111100100011110101001111000101",
    942 => "00111100011101011001100010011110",
    943 => "10111001011101111011110100100100",
    944 => "10101110010000101001011011111011",
    945 => "10111101111001011001010000010010",
    946 => "00111011110011101100000010000011",
    947 => "00110001001111010010111110101110",
    948 => "00111111011111100110001011101110",
    949 => "00111110000011101001010001101000",
    950 => "00111100100011110101001111000101",
    951 => "00111100011101011001100010011110",
    952 => "00111111011001110001101100100000",
    953 => "00111110011001000111111000110010",
    954 => "00111000111111110101110100010011",
    955 => "00111111011001110001101100100000",
    956 => "00111101010010111000010111101011",
    957 => "00110111010000110011111101100101",
    958 => "00111110000011101001010001101000",
    959 => "00111100100011110101001111000101",
    960 => "00111100011101011001100010011110",
    961 => "10111001011101111011101111010000",
    962 => "10101110010000101001010010001000",
    963 => "10111101111001011001001110101001",
    964 => "00111011110011101011111111000100",
    965 => "00110001001111010010110110100011",
    966 => "00111111011111100110001011101111",
    967 => "00111110000011101001010001101000",
    968 => "00111100100011110101001111000101",
    969 => "00111100011101011001100010011110",
    970 => "00111111011001110001101100011001",
    971 => "00111110011001000111111001000101",
    972 => "00111000111111110101110101001111",
    973 => "00111111011001110001101100011001",
    974 => "00111101010010111000011000000101",
    975 => "00110111010000110011111110011101",
    976 => "00111110000011101001010001101000",
    977 => "00111100100011110101001111000101",
    978 => "00111100011101011001100010011110",
    979 => "10111001011101111011101111010000",
    980 => "10101110010000101001010010001000",
    981 => "10111101111001011001001110101001",
    982 => "00111011110011101011111111000100",
    983 => "00110001001111010010110110100011",
    984 => "00111111011111100110001011101111",
    985 => "00111110000011101001010001101000",
    986 => "00111100100011110101001111000101",
    987 => "00111100011101011001100010011110",
    988 => "00111111011001110001101100011001",
    989 => "00111110011001000111111001000101",
    990 => "00111000111111110101110101001111",
    991 => "00111111011001110001101100011001",
    992 => "00111101010010111000011000000101",
    993 => "00110111010000110011111110011101",
    994 => "00111110110000001110110111111010",
    995 => "10111101010111000110010001101001",
    996 => "00111111011011001011101010111100",
    997 => "00111110000011101001010001101000",
    998 => "00111100100011110101001111000101",
    999 => "00111100011101011001100010011110");

  constant ans_lut : lut := (
    0 => "00111111011100000110011101110100",
    1 => "00111111011100001000111111010100",
    2 => "00111110101011110001011011100111",
    3 => "00111110101011110001110010001100",
    4 => "00111111010111001110100011000100",
    5 => "00111111010111011011010000100000",
    6 => "00111110111111111101010001001100",
    7 => "00111110111111111111111100000000",
    8 => "10111110111111111111111100000000",
    9 => "10111110101011110001110010001100",
    10 => "10111111011100001000111111010100",
    11 => "11000011001000111111011111010000",
    12 => "01000010110011101100111001001101",
    13 => "11000011001101101100001010111101",
    14 => "00111111001100101011100110110010",
    15 => "00111111010000011001110010011110",
    16 => "00111111010001000001101011100100",
    17 => "10111111010001000001101011100100",
    18 => "00111111001100101011100110110010",
    19 => "00111111001001000011010011100111",
    20 => "00111111001001001000111001110000",
    21 => "00111111001100101011100110110010",
    22 => "00111111010000011001110010011110",
    23 => "00111111010001000001101011100100",
    24 => "00111111001100101011100110110010",
    25 => "00111111001001000011010011100111",
    26 => "00111111001001001000111001110000",
    27 => "10111111000011100000000011010110",
    28 => "10111111100000000000000000000000",
    29 => "00111111011001100110011001101000",
    30 => "10111101001110100000110100100110",
    31 => "10111110001001010000000010100000",
    32 => "00111111101001111000110101110011",
    33 => "10111110000001011010100011000011",
    34 => "10111110000001011010100011011000",
    35 => "00111110000001011010100011011000",
    36 => "00111111011111011100111010000110",
    37 => "00111111011111011100111101010011",
    38 => "10111111011111011100111101010011",
    39 => "10111101001111010101011011000010",
    40 => "10111110001001100101001000100100",
    41 => "00111111101001100011101101110000",
    42 => "00111110110011011100111111001000",
    43 => "00111111011010110101000100110010",
    44 => "00111111011010111001100000011100",
    45 => "00111110110011011100111111001000",
    46 => "00111110110010000100010011011011",
    47 => "00111110110010000101000001000111",
    48 => "10111101110100101000100100000100",
    49 => "10111110000100110011010100101010",
    50 => "00111111011010001000000110101110",
    51 => "10111101101110011011111111100001",
    52 => "10111101101110011011111111101000",
    53 => "00111101101110011011111111101000",
    54 => "00111111011111101111000110110100",
    55 => "00111111011111101111000111100100",
    56 => "10111111011111101111000111100100",
    57 => "10111101010001000011001011110000",
    58 => "10111110001010001110110111000100",
    59 => "00111111101000111011101001011000",
    60 => "00111110110101101101001110111000",
    61 => "00111111011010010111011100101011",
    62 => "00111111011010011100101101001110",
    63 => "00111110110101101101001110111000",
    64 => "00111110110100001000011000001011",
    65 => "00111110110100001001010000110000",
    66 => "10111101110100001001111110000100",
    67 => "10111110000101010101000011110010",
    68 => "00111111011011000100010001011010",
    69 => "10111101101111001011111011001010",
    70 => "10111101101111001011111011010001",
    71 => "00111101101111001011111011010001",
    72 => "00111111011111101110100011100100",
    73 => "00111111011111101110100100010110",
    74 => "10111111011111101110100100010110",
    75 => "10111101010001000000010110010000",
    76 => "10111110001010001101110100100100",
    77 => "00111111101000111100100111011101",
    78 => "00111110110101101001101111011100",
    79 => "00111111011010011000001011100010",
    80 => "00111111011010011101011010101110",
    81 => "00111110110101101001101111011100",
    82 => "00111110110100000101001100011000",
    83 => "00111110110100000110000100101011",
    84 => "10111101110100001010101010011001",
    85 => "10111110000101010100010011100110",
    86 => "00111111011011000010111011110000",
    87 => "10111101101111001010110110111010",
    88 => "10111101101111001010110111000001",
    89 => "00111101101111001010110111000001",
    90 => "00111111011111101110100100010110",
    91 => "00111111011111101110100101001000",
    92 => "10111111011111101110100101001000",
    93 => "10111101010001000000011010011010",
    94 => "10111110001010001101110110000100",
    95 => "00111111101000111100100110000101",
    96 => "00111110110101101001110100011000",
    97 => "00111111011010011000001010100000",
    98 => "00111111011010011101011001101110",
    99 => "00111110110101101001110100011000",
    100 => "00111110110100000101010000111000",
    101 => "00111110110100000110001001001011",
    102 => "10111101110100001010101001011010",
    103 => "10111110000101010100010100101010",
    104 => "00111111011011000010111101101010",
    105 => "10111101101111001010111000011100",
    106 => "10111101101111001010111000100011",
    107 => "00111101101111001010111000100011",
    108 => "00111111011111101110100100010101",
    109 => "00111111011111101110100101001000",
    110 => "10111111011111101110100101001000",
    111 => "10111101010001000000011010010010",
    112 => "10111110001010001101110110000010",
    113 => "00111111101000111100100110000110",
    114 => "00111110110101101001110100010100",
    115 => "00111111011010011000001010100000",
    116 => "00111111011010011101011001101110",
    117 => "00111110110101101001110100010100",
    118 => "00111110110100000101010000110101",
    119 => "00111110110100000110001001001000",
    120 => "10111111000101100111110100111110",
    121 => "00111101011100101101101011101100",
    122 => "10111111010011101000101000101010",
    123 => "10111101001110100000110100100110",
    124 => "10111110001001010000000010100000",
    125 => "00111111101001111000110101110011",
    126 => "00111110110010010000111011111000",
    127 => "00111111011011000100001011110000",
    128 => "00111111011011001000001110001010",
    129 => "00111110110010010000111011111000",
    130 => "00111110110000111110010000011010",
    131 => "00111110110000111110111001000100",
    132 => "10111101110100111010001001011110",
    133 => "10111110000100011111011111110010",
    134 => "00111111011001100100100011111000",
    135 => "00111111010000101101111000000011",
    136 => "00111111001101011101010101100001",
    137 => "00111111001110010101100010100010",
    138 => "00111111010000101101111000000011",
    139 => "00111111001100000000110001110110",
    140 => "00111111001100001001011000011111",
    141 => "10111101110110110101100011001100",
    142 => "10111110000010001011011010010111",
    143 => "00111111010101010111010101101100",
    144 => "00111111001011100001010010111110",
    145 => "00111111001011101001010011111111",
    146 => "00111111001101111110101001010110",
    147 => "00111111001110110011110001000111",
    148 => "10111101110110101110011111110010",
    149 => "10111110000010010100010011000010",
    150 => "00111111010101100111101010000110",
    151 => "00111111001011101011110101000000",
    152 => "00111111001011110100000010010100",
    153 => "00111111001101110011100110010000",
    154 => "00111111001110101001101110110110",
    155 => "10111101110110101110111110010110",
    156 => "10111110000010010011101100101010",
    157 => "00111111010101100110100011101010",
    158 => "00111111001011101011000111100111",
    159 => "00111111001011110011010100000110",
    160 => "00111111001101110100010110000100",
    161 => "00111111001110101010011010010000",
    162 => "10111101110110101110111100010100",
    163 => "10111110000010010011101111001100",
    164 => "00111111010101100110101000010100",
    165 => "00111111001011101011001010101000",
    166 => "00111111001011110011010111001010",
    167 => "00111111001101110100010010111000",
    168 => "00111111001110101010010111010110",
    169 => "10111101110110101110111100011101",
    170 => "10111110000010010011101111000010",
    171 => "00111111010101100110101000000000",
    172 => "00111111001011101011001010011010",
    173 => "00111111001011110011010110111100",
    174 => "00111111001101110100010011000110",
    175 => "00111111001110101010010111100011",
    176 => "10111101110110101110111100011100",
    177 => "10111110000010010011101111000011",
    178 => "00111111010101100110101000000010",
    179 => "00111111001011101011001010011101",
    180 => "00111111001011110011010110111111",
    181 => "00111111001101110100010011000100",
    182 => "00111111001110101010010111100001",
    183 => "10111101110110101110111100011101",
    184 => "10111110000010010011101111000010",
    185 => "00111111010101100110101000000000",
    186 => "00111111001011101011001010011010",
    187 => "00111111001011110011010110111100",
    188 => "00111111001101110100010011000110",
    189 => "00111111001110101010010111100011",
    190 => "10111101110110101110111100011100",
    191 => "10111110000010010011101111000011",
    192 => "00111111010101100110101000000010",
    193 => "00111111001011101011001010011101",
    194 => "00111111001011110011010110111111",
    195 => "00111111001101110100010011000100",
    196 => "00111111001110101010010111100001",
    197 => "10111111000010111110011110000001",
    198 => "10111111000010111110011101111111",
    199 => "10111111001000100111001011100000",
    200 => "10111110100110011001100110011000",
    201 => "10111101001110100000110100100110",
    202 => "10111110001001010000000010100000",
    203 => "00111111101001111000110101110011",
    204 => "10111110110000111110010100101100",
    205 => "10111110110000111110111101010110",
    206 => "00111110110000111110111101010110",
    207 => "00111111011011000100001010110101",
    208 => "00111111011011001000001101010001",
    209 => "10111111011011001000001101010001",
    210 => "10111101010101110100110101100010",
    211 => "10111110001011110010101110101110",
    212 => "00111111100111100100111011110111",
    213 => "00111110111010100101011001001100",
    214 => "00111111011001010010111111000100",
    215 => "00111111011001011010011011000011",
    216 => "00111110111010100101011001001100",
    217 => "00111110111000100010011111010101",
    218 => "00111110111000100011110110101000",
    219 => "10111101110011011001001110011100",
    220 => "10111110000110001000110100100110",
    221 => "00111111011100011111110000101100",
    222 => "10111110100011110011111010111101",
    223 => "10111110100011110100000010111101",
    224 => "00111110100011110100000010111101",
    225 => "00111111011101011011010011110010",
    226 => "00111111011101011100011010001110",
    227 => "10111111011101011100011010001110",
    228 => "10111101100000000000010111010001",
    229 => "10111110001101110111011101110110",
    230 => "00111111100101111111100010100101",
    231 => "00111111000000001001001101010010",
    232 => "00111111010111111011011000101100",
    233 => "00111111011000000110001001111010",
    234 => "00111111000000001001001101010010",
    235 => "00111110111101100101011011111001",
    236 => "00111110111101100111100110101100",
    237 => "10111101110011100110111011111010",
    238 => "10111110000101111010100000101000",
    239 => "00111111011100000110100100011100",
    240 => "10111110100011100101011010001111",
    241 => "10111110100011100101100001111110",
    242 => "00111110100011100101100001111110",
    243 => "00111111011101011101011100100000",
    244 => "00111111011101011110100001001000",
    245 => "10111111011101011110100001001000",
    246 => "10111101100000000011101001011101",
    247 => "10111110001101111000001111110110",
    248 => "00111111100101111110110111111101",
    249 => "00111111000000001010011010000000",
    250 => "00111111010111111010110010001010",
    251 => "00111111011000000101100100111110",
    252 => "00111111000000001010011010000000",
    253 => "00111110111101100111100001111110",
    254 => "00111110111101101001101101001011",
    255 => "10111101110011100111100101000101",
    256 => "10111110000101111001110101010100",
    257 => "00111111011100000101011000000110",
    258 => "10111110100011100100101110010000",
    259 => "10111110100011100100110101111111",
    260 => "00111110100011100100110101111111",
    261 => "00111111011101011101100010111101",
    262 => "00111111011101011110100111100000",
    263 => "10111111011101011110100111100000",
    264 => "10111101100000000011110011010011",
    265 => "10111110001101111000010010001010",
    266 => "00111111100101111110110101111110",
    267 => "00111111000000001010011101100110",
    268 => "00111111010111111010110000010110",
    269 => "00111111011000000101100011001111",
    270 => "00111111000000001010011101100110",
    271 => "00111110111101100111101000010000",
    272 => "00111110111101101001110011011110",
    273 => "10111101110011100111100111000000",
    274 => "10111110000101111001110011010010",
    275 => "00111111011100000101010100100010",
    276 => "10111110100011100100101100001101",
    277 => "10111110100011100100110011111011",
    278 => "00111110100011100100110011111011",
    279 => "00111111011101011101100011010000",
    280 => "00111111011101011110100111110010",
    281 => "10111111011101011110100111110010",
    282 => "10111101100000000011110011110000",
    283 => "10111110001101111000010010010010",
    284 => "00111111100101111110110101111000",
    285 => "00111111000000001010011101110000",
    286 => "00111111010111111010110000010001",
    287 => "00111111011000000101100011001010",
    288 => "00111111000000001010011101110000",
    289 => "00111110111101100111101000100001",
    290 => "00111110111101101001110011101111",
    291 => "10111111000100010000100001100001",
    292 => "00111110001101111111110000110011",
    293 => "10111111010011011110000011010100",
    294 => "10111101001110100000110100100110",
    295 => "10111110001001010000000010100000",
    296 => "00111111101001111000110101110011",
    297 => "00111111001001111000110011011011",
    298 => "00111111010010010010101101110110",
    299 => "00111111010010110001100101101110",
    300 => "00111111001001111000110011011011",
    301 => "00111111000110111001011010010100",
    302 => "00111111000110111101011110000001",
    303 => "10111101101010000011001001011000",
    304 => "10111110001100111100111101100110",
    305 => "00111111100011111000001100101100",
    306 => "00111111000011111100110100101100",
    307 => "00111111010101111001110010010010",
    308 => "00111111010110001010100110011010",
    309 => "00111111000011111100110100101100",
    310 => "00111111000010000011110100110011",
    311 => "00111111000010000101101110000100",
    312 => "10111101110110000110101110101101",
    313 => "10111110000011000101011100001110",
    314 => "00111111010111000001100011110100",
    315 => "00111111000100001100010010000110",
    316 => "00111111000100001110111101000110",
    317 => "00111111010100011010001101111101",
    318 => "00111111010100110000010101101110",
    319 => "10111101110001000110010111001100",
    320 => "10111110001000010110000000001100",
    321 => "00111111100000001001101100110100",
    322 => "00111111001010101010000111101010",
    323 => "00111111010001110010001001000111",
    324 => "00111111010010010011010101010100",
    325 => "00111111001010101010000111101010",
    326 => "00111111000111011111111110000010",
    327 => "00111111000111100100011010011010",
    328 => "10111101110110111000100100110100",
    329 => "10111110000010000111100101011010",
    330 => "00111111010101010000010011011100",
    331 => "00111111000011001010111001111000",
    332 => "00111111000011001101001011001011",
    333 => "00111111010101001001001010011100",
    334 => "00111111010101011100100101100111",
    335 => "10111101110001001011011110101011",
    336 => "10111110001000010001011101010010",
    337 => "00111111100000000101110110100100",
    338 => "00111111001010110001000010111011",
    339 => "00111111010001101101100001010010",
    340 => "00111111010010001111000010111110",
    341 => "00111111001010110001000010111011",
    342 => "00111111000111100101010110100101",
    343 => "00111111000111101001110110100100",
    344 => "10111101110110111000101100100110",
    345 => "10111110000010000111011011100010",
    346 => "00111111010101010000000001010010",
    347 => "00111111000011001010101111010101",
    348 => "00111111000011001101000000100011",
    349 => "00111111010101001001010001110110",
    350 => "00111111010101011100101100100111",
    351 => "10111101110001001011011111011000",
    352 => "10111110001000010001011100101000",
    353 => "00111111100000000101110110000011",
    354 => "00111111001010110001000011110110",
    355 => "00111111010001101101100000101011",
    356 => "00111111010010001111000010011010",
    357 => "00111111001010110001000011110110",
    358 => "00111111000111100101010111010011",
    359 => "00111111000111101001110111010010",
    360 => "10111101110110111000101100101000",
    361 => "10111110000010000111011011100000",
    362 => "00111111010101010000000001001110",
    363 => "00111111000011001010101111010011",
    364 => "00111111000011001101000000100001",
    365 => "00111111010101001001010001111000",
    366 => "00111111010101011100101100101001",
    367 => "10111101110001001011011111011011",
    368 => "10111110001000010001011100100110",
    369 => "00111111100000000101110110000001",
    370 => "00111111001010110001000011111010",
    371 => "00111111010001101101100000101000",
    372 => "00111111010010001111000010010110",
    373 => "00111111001010110001000011111010",
    374 => "00111111000111100101010111010110",
    375 => "00111111000111101001110111010101",
    376 => "10111111000110001010111000000001",
    377 => "10111110110101011111110011001000",
    378 => "10111111001011110110111100111100",
    379 => "10111110111111111111111111111110",
    380 => "10111101001110100000110100100110",
    381 => "10111110001001010000000010100000",
    382 => "00111111101001111000110101110011",
    383 => "10111111000110111001011100001010",
    384 => "10111111000110111101011111111000",
    385 => "00111111000110111101011111111000",
    386 => "00111111010010010010101100010100",
    387 => "00111111010010110001100100010011",
    388 => "10111111010010110001100100010011",
    389 => "10111101100001001011101011011000",
    390 => "10111110001110000110100101111110",
    391 => "00111111100101110001001100110100",
    392 => "00111111000000100011000001010010",
    393 => "00111111010111101110010101110010",
    394 => "00111111010111111001101010000110",
    395 => "00111111000000100011000001010010",
    396 => "00111110111110010010011101111011",
    397 => "00111110111110010100110001101000",
    398 => "10111101110011110111001010001000",
    399 => "10111110000101101001010100110100",
    400 => "00111111011011101000001101110010",
    401 => "10111110111001011110001011111100",
    402 => "10111110111001011111101011010011",
    403 => "00111110111001011111101011010011",
    404 => "00111111011001000011100011101011",
    405 => "00111111011001001011100010010111",
    406 => "10111111011001001011100010010111",
    407 => "10111101101001001011100100101000",
    408 => "10111110001101010010110011100010",
    409 => "00111111100100001001110100011100",
    410 => "00111111000011011101000110110000",
    411 => "00111111010110001011011110101100",
    412 => "00111111010110011011011000111111",
    413 => "00111111000011011101000110110000",
    414 => "00111111000001101001000010101110",
    415 => "00111111000001101010110011110111",
    416 => "10111101110101111011001010000110",
    417 => "10111110000011010011011011111010",
    418 => "00111111010111011011000010111110",
    419 => "10111110110101101100001101100111",
    420 => "10111110110101101101001111110011",
    421 => "00111110110101101101001111110011",
    422 => "00111111011010000000000010101100",
    423 => "00111111011010000110000000001110",
    424 => "10111111011010000110000000001110",
    425 => "10111101101001101100101010110000",
    426 => "10111110001101000110001011100010",
    427 => "00111111100011111111100100110010",
    428 => "00111111000011101111100010111010",
    429 => "00111111010110000001001110010000",
    430 => "00111111010110010001101001111000",
    431 => "00111111000011101111100010111010",
    432 => "00111111000001111000101000010100",
    433 => "00111111000001111010011110001000",
    434 => "10111101110110000010001011011101",
    435 => "10111110000011001010111101100000",
    436 => "00111111010111001011100111101000",
    437 => "10111110110101011110001110011011",
    438 => "10111110110101011111001111001100",
    439 => "00111110110101011111001111001100",
    440 => "00111111011010000011010111111111",
    441 => "00111111011010001001001110111100",
    442 => "10111111011010001001001110111100",
    443 => "10111101101001101110010010111011",
    444 => "10111110001101000101100001111010",
    445 => "00111111100011111111000011010111",
    446 => "00111111000011110000011111000110",
    447 => "00111111010110000000101100101000",
    448 => "00111111010110010001001001111111",
    449 => "00111111000011110000011111000110",
    450 => "00111111000001111001011011000111",
    451 => "00111111000001111011010001001010",
    452 => "10111101110110000010100000111111",
    453 => "10111110000011001010100011011011",
    454 => "00111111010111001010111000001000",
    455 => "10111110110101011101100011010101",
    456 => "10111110110101011110100100000010",
    457 => "00111110110101011110100100000010",
    458 => "00111111011010000011100010001110",
    459 => "00111111011010001001011000110111",
    460 => "10111111011010001001011000110111",
    461 => "10111101101001101110010111111000",
    462 => "10111110001101000101011111111100",
    463 => "00111111100011111111000001110001",
    464 => "00111111000011110000100001111100",
    465 => "00111111010110000000101011000010",
    466 => "00111111010110010001001000011110",
    467 => "00111111000011110000100001111100",
    468 => "00111111000001111001011101100000",
    469 => "00111111000001111011010011100100",
    470 => "10111111000110110001111110000110",
    471 => "00111110100110001101110011011001",
    472 => "10111111001111001100001100010000",
    473 => "10111101001110100000110100100110",
    474 => "10111110001001010000000010100000",
    475 => "00111111101001111000110101110011",
    476 => "00111111000110111001011100001100",
    477 => "00111111000110111101011111111010",
    478 => "00111111010010010010101100010010",
    479 => "00111111010010110001100100010001",
    480 => "10111101100001001011101011011000",
    481 => "10111110001110000110100101111110",
    482 => "00111111100101110001001100110100",
    483 => "00111111000000100011000001010010",
    484 => "00111111010111101110010101110010",
    485 => "00111111010111111001101010000110",
    486 => "00111111000000100011000001010010",
    487 => "00111110111110010010011101111011",
    488 => "00111110111110010100110001101000",
    489 => "10111101110011110111001010001000",
    490 => "10111110000101101001010100110100",
    491 => "00111111011011101000001101110010",
    492 => "00111110111001011110001011111111",
    493 => "00111110111001011111101011010110",
    494 => "00111111011001000011100011101010",
    495 => "00111111011001001011100010010110",
    496 => "10111101101001001011100100101010",
    497 => "10111110001101010010110011100010",
    498 => "00111111100100001001110100011011",
    499 => "00111111000011011101000110110010",
    500 => "00111111010110001011011110101011",
    501 => "00111111010110011011011000111110",
    502 => "00111111000011011101000110110010",
    503 => "00111111000001101001000010110000",
    504 => "00111111000001101010110011111001",
    505 => "10111101110101111011001010000110",
    506 => "10111110000011010011011011111010",
    507 => "00111111010111011011000010111110",
    508 => "00111110110101101100001101101010",
    509 => "00111110110101101101001111110110",
    510 => "00111111011010000000000010101100",
    511 => "00111111011010000110000000001110",
    512 => "10111101101001101100101010110001",
    513 => "10111110001101000110001011100000",
    514 => "00111111100011111111100100110011",
    515 => "00111111000011101111100010111000",
    516 => "00111111010110000001001110010001",
    517 => "00111111010110010001101001111000",
    518 => "00111111000011101111100010111000",
    519 => "00111111000001111000101000010010",
    520 => "00111111000001111010011110000110",
    521 => "10111101110110000010001011011110",
    522 => "10111110000011001010111101011111",
    523 => "00111111010111001011100111100110",
    524 => "00111110110101011110001110011100",
    525 => "00111110110101011111001111001110",
    526 => "00111111011010000011010111111110",
    527 => "00111111011010001001001110111010",
    528 => "10111101101001101110010010111110",
    529 => "10111110001101000101100001111010",
    530 => "00111111100011111111000011010101",
    531 => "00111111000011110000011111001000",
    532 => "00111111010110000000101100100111",
    533 => "00111111010110010001001001111101",
    534 => "00111111000011110000011111001000",
    535 => "00111111000001111001011011001000",
    536 => "00111111000001111011010001001011",
    537 => "10111101110110000010100000111111",
    538 => "10111110000011001010100011011011",
    539 => "00111111010111001010111000001000",
    540 => "00111110110101011101100011011000",
    541 => "00111110110101011110100100000101",
    542 => "00111111011010000011100010001101",
    543 => "00111111011010001001011000110110",
    544 => "10111101101001101110010111111010",
    545 => "10111110001101000101011111111010",
    546 => "00111111100011111111000001110001",
    547 => "00111111000011110000100001111100",
    548 => "00111111010110000000101011000010",
    549 => "00111111010110010001001000011110",
    550 => "00111111000011110000100001111100",
    551 => "00111111000001111001011101100000",
    552 => "00111111000001111011010011100100",
    553 => "10111111000110110001111110001000",
    554 => "10111110100110001101110011011100",
    555 => "10111111001111001100001100010000",
    556 => "10111111001100110011001100110010",
    557 => "10111101001110100000110100100110",
    558 => "10111110001001010000000010100000",
    559 => "00111111101001111000110101110011",
    560 => "10111111010010011011111110010110",
    561 => "10111111010010110001100101100000",
    562 => "00111111010010110001100101100000",
    563 => "00111111000101001000011110100000",
    564 => "00111111000110111101011101010110",
    565 => "10111111000110111101011101010110",
    566 => "10111101101010000011001001100111",
    567 => "10111110001100111100111101100000",
    568 => "00111111100011111000001100101000",
    569 => "00111111000011111100110100110100",
    570 => "00111111010101111001110010001110",
    571 => "00111111010110001010100110010110",
    572 => "00111111000011111100110100110100",
    573 => "00111111000010000011110100111010",
    574 => "00111111000010000101101110001011",
    575 => "10111101110110000110101110110001",
    576 => "10111110000011000101011100001001",
    577 => "00111111010111000001100011101110",
    578 => "10111111000100001100010010000010",
    579 => "10111111000100001110111101000010",
    580 => "00111111000100001110111101000010",
    581 => "00111111010100011010001110000000",
    582 => "00111111010100110000010101110000",
    583 => "10111111010100110000010101110000",
    584 => "10111101110001000110010111001110",
    585 => "10111110001000010110000000001100",
    586 => "00111111100000001001101100110011",
    587 => "00111111001010101010000111101100",
    588 => "00111111010001110010001001000110",
    589 => "00111111010010010011010101010010",
    590 => "00111111001010101010000111101100",
    591 => "00111111000111011111111110000011",
    592 => "00111111000111100100011010011011",
    593 => "10111101110110111000100100110100",
    594 => "10111110000010000111100101011010",
    595 => "00111111010101010000010011011100",
    596 => "10111111000011001010111001110111",
    597 => "10111111000011001101001011001001",
    598 => "00111111000011001101001011001001",
    599 => "00111111010101001001001010011110",
    600 => "00111111010101011100100101101001",
    601 => "10111111010101011100100101101001",
    602 => "10111101110001001011011110101001",
    603 => "10111110001000010001011101010010",
    604 => "00111111100000000101110110100110",
    605 => "00111111001010110001000010110111",
    606 => "00111111010001101101100001010101",
    607 => "00111111010010001111000011000001",
    608 => "00111111001010110001000010110111",
    609 => "00111111000111100101010110100010",
    610 => "00111111000111101001110110100000",
    611 => "10111101110110111000101100100110",
    612 => "10111110000010000111011011100010",
    613 => "00111111010101010000000001010010",
    614 => "10111111000011001010101111010100",
    615 => "10111111000011001101000000100011",
    616 => "00111111000011001101000000100011",
    617 => "00111111010101001001010001110111",
    618 => "00111111010101011100101100101000",
    619 => "10111111010101011100101100101000",
    620 => "10111101110001001011011111011010",
    621 => "10111110001000010001011100101000",
    622 => "00111111100000000101110110000001",
    623 => "00111111001010110001000011111010",
    624 => "00111111010001101101100000101000",
    625 => "00111111010010001111000010010110",
    626 => "00111111001010110001000011111010",
    627 => "00111111000111100101010111010110",
    628 => "00111111000111101001110111010101",
    629 => "10111101110110111000101100100110",
    630 => "10111110000010000111011011100010",
    631 => "00111111010101010000000001010010",
    632 => "10111111000011001010101111010100",
    633 => "10111111000011001101000000100011",
    634 => "00111111000011001101000000100011",
    635 => "00111111010101001001010001110111",
    636 => "00111111010101011100101100101000",
    637 => "10111111010101011100101100101000",
    638 => "10111101110001001011011111011010",
    639 => "10111110001000010001011100101000",
    640 => "00111111100000000101110110000001",
    641 => "00111111001010110001000011111010",
    642 => "00111111010001101101100000101000",
    643 => "00111111010010001111000010010110",
    644 => "00111111001010110001000011111010",
    645 => "00111111000111100101010111010110",
    646 => "00111111000111101001110111010101",
    647 => "10111111000110001010111000000001",
    648 => "00111110110101011111110011000110",
    649 => "10111111001011110110111100111110",
    650 => "10111101001110100000110100100110",
    651 => "10111110001001010000000010100000",
    652 => "00111111101001111000110101110011",
    653 => "00111110110000111110010100101110",
    654 => "00111110110000111110111101011000",
    655 => "00111111011011000100001010110101",
    656 => "00111111011011001000001101010001",
    657 => "10111101010101110100110101100010",
    658 => "10111110001011110010101110101110",
    659 => "00111111100111100100111011110111",
    660 => "00111110111010100101011001001100",
    661 => "00111111011001010010111111000100",
    662 => "00111111011001011010011011000011",
    663 => "00111110111010100101011001001100",
    664 => "00111110111000100010011111010101",
    665 => "00111110111000100011110110101000",
    666 => "10111101110011011001001110011100",
    667 => "10111110000110001000110100100110",
    668 => "00111111011100011111110000101100",
    669 => "00111110100011110011111010111111",
    670 => "00111110100011110100000010111111",
    671 => "00111111011101011011010011110010",
    672 => "00111111011101011100011010001110",
    673 => "10111101100000000000010111010011",
    674 => "10111110001101110111011101110110",
    675 => "00111111100101111111100010100101",
    676 => "00111111000000001001001101010010",
    677 => "00111111010111111011011000101100",
    678 => "00111111011000000110001001111010",
    679 => "00111111000000001001001101010010",
    680 => "00111110111101100101011011111001",
    681 => "00111110111101100111100110101100",
    682 => "10111101110011100110111011111010",
    683 => "10111110000101111010100000101000",
    684 => "00111111011100000110100100011100",
    685 => "00111110100011100101011010010001",
    686 => "00111110100011100101100010000000",
    687 => "00111111011101011101011100100000",
    688 => "00111111011101011110100001001000",
    689 => "10111101100000000011101001011111",
    690 => "10111110001101111000001111110110",
    691 => "00111111100101111110110111111101",
    692 => "00111111000000001010011010000000",
    693 => "00111111010111111010110010001010",
    694 => "00111111011000000101100100111110",
    695 => "00111111000000001010011010000000",
    696 => "00111110111101100111100001111110",
    697 => "00111110111101101001101101001011",
    698 => "10111101110011100111100101000101",
    699 => "10111110000101111001110101010100",
    700 => "00111111011100000101011000000110",
    701 => "00111110100011100100101110010010",
    702 => "00111110100011100100110110000001",
    703 => "00111111011101011101100010111101",
    704 => "00111111011101011110100111100000",
    705 => "10111101100000000011110011010011",
    706 => "10111110001101111000010010001010",
    707 => "00111111100101111110110101111110",
    708 => "00111111000000001010011101100110",
    709 => "00111111010111111010110000010110",
    710 => "00111111011000000101100011001111",
    711 => "00111111000000001010011101100110",
    712 => "00111110111101100111101000010000",
    713 => "00111110111101101001110011011110",
    714 => "10111101110011100111100111000000",
    715 => "10111110000101111001110011010010",
    716 => "00111111011100000101010100100010",
    717 => "00111110100011100100101100001111",
    718 => "00111110100011100100110011111101",
    719 => "00111111011101011101100011010000",
    720 => "00111111011101011110100111110010",
    721 => "10111101100000000011110011110010",
    722 => "10111110001101111000010010010010",
    723 => "00111111100101111110110101110111",
    724 => "00111111000000001010011101110010",
    725 => "00111111010111111010110000010000",
    726 => "00111111011000000101100011001010",
    727 => "00111111000000001010011101110010",
    728 => "00111110111101100111101000100100",
    729 => "00111110111101101001110011110010",
    730 => "10111111000100010000100001100010",
    731 => "10111110001101111111110000110110",
    732 => "10111111010011011110000011010100",
    733 => "10111111011001100110011001100110",
    734 => "10111101001110100000110100100110",
    735 => "10111110001001010000000010100000",
    736 => "00111111101001111000110101110011",
    737 => "10111111011001111101010001000010",
    738 => "10111111011011001000001100101001",
    739 => "00111111011011001000001100101001",
    740 => "00111110100111001011000010111000",
    741 => "00111110110000111110100001011100",
    742 => "10111110110000111110100001011100",
    743 => "10111101110100111010010000101000",
    744 => "10111110000100011111010111101010",
    745 => "00111111011001100100010101010010",
    746 => "00111111010000101110000101001011",
    747 => "00111111001101011101001011100010",
    748 => "00111111001110010101011001011111",
    749 => "00111111010000101110000101001011",
    750 => "00111111001100000000111011001011",
    751 => "00111111001100001001100010000000",
    752 => "10111101110110110101100010111000",
    753 => "10111110000010001011011010110000",
    754 => "00111111010101010111010110011010",
    755 => "10111111001011100001010011011100",
    756 => "10111111001011101001010100011101",
    757 => "00111111001011101001010100011101",
    758 => "00111111001101111110101000110110",
    759 => "00111111001110110011110000101010",
    760 => "10111111001110110011110000101010",
    761 => "10111101110110101110011111110100",
    762 => "10111110000010010100010011000010",
    763 => "00111111010101100111101010000100",
    764 => "00111111001011101011110100111111",
    765 => "00111111001011110100000010010011",
    766 => "00111111001101110011100110010010",
    767 => "00111111001110101001101110111000",
    768 => "10111101110110101110111110010110",
    769 => "10111110000010010011101100101010",
    770 => "00111111010101100110100011101010",
    771 => "10111111001011101011000111100111",
    772 => "10111111001011110011010100000110",
    773 => "00111111001011110011010100000110",
    774 => "00111111001101110100010110000100",
    775 => "00111111001110101010011010010000",
    776 => "10111111001110101010011010010000",
    777 => "10111101110110101110111100010100",
    778 => "10111110000010010011101111001110",
    779 => "00111111010101100110101000010110",
    780 => "00111111001011101011001010101010",
    781 => "00111111001011110011010111001100",
    782 => "00111111001101110100010010110110",
    783 => "00111111001110101010010111010100",
    784 => "10111101110110101110111100011111",
    785 => "10111110000010010011101111000000",
    786 => "00111111010101100110100111111010",
    787 => "10111111001011101011001010010110",
    788 => "10111111001011110011010110111000",
    789 => "00111111001011110011010110111000",
    790 => "00111111001101110100010011001011",
    791 => "00111111001110101010010111100111",
    792 => "10111111001110101010010111100111",
    793 => "10111101110110101110111100011011",
    794 => "10111110000010010011101111000100",
    795 => "00111111010101100110101000000100",
    796 => "00111111001011101011001010011110",
    797 => "00111111001011110011010111000000",
    798 => "00111111001101110100010011000011",
    799 => "00111111001110101010010111100000",
    800 => "10111101110110101110111100011100",
    801 => "10111110000010010011101111000011",
    802 => "00111111010101100110101000000010",
    803 => "10111111001011101011001010011011",
    804 => "10111111001011110011010110111101",
    805 => "00111111001011110011010110111101",
    806 => "00111111001101110100010011000110",
    807 => "00111111001110101010010111100011",
    808 => "10111111001110101010010111100011",
    809 => "10111101110110101110111100011100",
    810 => "10111110000010010011101111000011",
    811 => "00111111010101100110101000000010",
    812 => "00111111001011101011001010011101",
    813 => "00111111001011110011010110111111",
    814 => "00111111001101110100010011000100",
    815 => "00111111001110101010010111100001",
    816 => "10111111000010111110011110000001",
    817 => "00111111000010111110011101111110",
    818 => "10111111001000100111001011100000",
    819 => "10111101001110100000110100100110",
    820 => "10111110001001010000000010100000",
    821 => "00111111101001111000110101110011",
    822 => "00111110000001011010100011000011",
    823 => "00111110000001011010100011011000",
    824 => "00111111011111011100111010000110",
    825 => "00111111011111011100111101010011",
    826 => "10111101001111010101011011000010",
    827 => "10111110001001100101001000100100",
    828 => "00111111101001100011101101110000",
    829 => "00111110110011011100111111001000",
    830 => "00111111011010110101000100110010",
    831 => "00111111011010111001100000011100",
    832 => "00111110110011011100111111001000",
    833 => "00111110110010000100010011011011",
    834 => "00111110110010000101000001000111",
    835 => "10111101110100101000100100000100",
    836 => "10111110000100110011010100101010",
    837 => "00111111011010001000000110101110",
    838 => "00111101101110011011111111100001",
    839 => "00111101101110011011111111101000",
    840 => "00111111011111101111000110110100",
    841 => "00111111011111101111000111100100",
    842 => "10111101010001000011001011110000",
    843 => "10111110001010001110110111000100",
    844 => "00111111101000111011101001011000",
    845 => "00111110110101101101001110111000",
    846 => "00111111011010010111011100101011",
    847 => "00111111011010011100101101001110",
    848 => "00111110110101101101001110111000",
    849 => "00111110110100001000011000001011",
    850 => "00111110110100001001010000110000",
    851 => "10111101110100001001111110000100",
    852 => "10111110000101010101000011110010",
    853 => "00111111011011000100010001011010",
    854 => "00111101101111001011111011001010",
    855 => "00111101101111001011111011010001",
    856 => "00111111011111101110100011100100",
    857 => "00111111011111101110100100010110",
    858 => "10111101010001000000010110010000",
    859 => "10111110001010001101110100100100",
    860 => "00111111101000111100100111011101",
    861 => "00111110110101101001101111011100",
    862 => "00111111011010011000001011100010",
    863 => "00111111011010011101011010101110",
    864 => "00111110110101101001101111011100",
    865 => "00111110110100000101001100011000",
    866 => "00111110110100000110000100101011",
    867 => "10111101110100001010101010011001",
    868 => "10111110000101010100010011100110",
    869 => "00111111011011000010111011110000",
    870 => "00111101101111001010110110111010",
    871 => "00111101101111001010110111000001",
    872 => "00111111011111101110100100010110",
    873 => "00111111011111101110100101001000",
    874 => "10111101010001000000011010011010",
    875 => "10111110001010001101110110000100",
    876 => "00111111101000111100100110000101",
    877 => "00111110110101101001110100011000",
    878 => "00111111011010011000001010100000",
    879 => "00111111011010011101011001101110",
    880 => "00111110110101101001110100011000",
    881 => "00111110110100000101010000111000",
    882 => "00111110110100000110001001001011",
    883 => "10111101110100001010101001011010",
    884 => "10111110000101010100010100101010",
    885 => "00111111011011000010111101101010",
    886 => "00111101101111001010111000011100",
    887 => "00111101101111001010111000100011",
    888 => "00111111011111101110100100010101",
    889 => "00111111011111101110100101001000",
    890 => "10111101010001000000011010010010",
    891 => "10111110001010001101110110000010",
    892 => "00111111101000111100100110000110",
    893 => "00111110110101101001110100010100",
    894 => "00111111011010011000001010100000",
    895 => "00111111011010011101011001101110",
    896 => "00111110110101101001110100010100",
    897 => "00111110110100000101010000110101",
    898 => "00111110110100000110001001001000",
    899 => "10111111000101100111110100111110",
    900 => "10111101011100101101101011101100",
    901 => "10111111010011101000101000101010",
    902 => "00111111001100110011001100110110",
    903 => "10111101110011001100110011000000",
    904 => "10111101001110100000110100100110",
    905 => "10111110001001010000000010100000",
    906 => "00111111101001111000110101110011",
    907 => "10111110000001011010100010111011",
    908 => "10111110000001011010100011010000",
    909 => "00111110000001011010100011010000",
    910 => "00111111011111011100111010000110",
    911 => "00111111011111011100111101010011",
    912 => "10111111011111011100111101010011",
    913 => "10111101001111010101011011000010",
    914 => "10111110001001100101001000100100",
    915 => "00111111101001100011101101110000",
    916 => "00111111001010010110011000010000",
    917 => "00111111010001111111010000001011",
    918 => "00111111010010011111100000000010",
    919 => "00111111001010010110011000010000",
    920 => "00111111000111010000100101010000",
    921 => "00111111000111010100110111100001",
    922 => "10111101101001111011101100011001",
    923 => "10111110001101000000000100111000",
    924 => "00111111100011111010101011101100",
    925 => "10111101111001010110001010101010",
    926 => "10111101111001010110001010111110",
    927 => "00111101111001010110001010111110",
    928 => "00111111011111100110001100110010",
    929 => "00111111011111100110001110100001",
    930 => "10111111011111100110001110100001",
    931 => "10111101010000000110110010001010",
    932 => "10111110001001111000010010000100",
    933 => "00111111101001010001000010110010",
    934 => "00111111001010110000100001001100",
    935 => "00111111010001101101110111110101",
    936 => "00111111010010001111010111111000",
    937 => "00111111001010110000100001001100",
    938 => "00111111000111100100111100011000",
    939 => "00111111000111101001011100000101",
    940 => "10111101101001110101110010111000",
    941 => "10111110001101000010100000000000",
    942 => "00111111100011111100100111110011",
    943 => "10111101111001011001001111111110",
    944 => "10111101111001011001010000010010",
    945 => "00111101111001011001010000010010",
    946 => "00111111011111100110001001111111",
    947 => "00111111011111100110001011101110",
    948 => "10111111011111100110001011101110",
    949 => "10111101010000000110010101001000",
    950 => "10111110001001111000000110111110",
    951 => "00111111101001010001001101011101",
    952 => "00111111001010110000010010010000",
    953 => "00111111010001101110000001110100",
    954 => "00111111010010001111100001001000",
    955 => "00111111001010110000010010010000",
    956 => "00111111000111100100110000110001",
    957 => "00111111000111101001010000010111",
    958 => "10111101101001110101110110000100",
    959 => "10111110001101000010011110101100",
    960 => "00111111100011111100100110110001",
    961 => "10111101111001011001001110010101",
    962 => "10111101111001011001001110101001",
    963 => "00111101111001011001001110101001",
    964 => "00111111011111100110001010000000",
    965 => "00111111011111100110001011101111",
    966 => "10111111011111100110001011101111",
    967 => "10111101010000000110010101011000",
    968 => "10111110001001111000000111000100",
    969 => "00111111101001010001001101011000",
    970 => "00111111001010110000010010010111",
    971 => "00111111010001101110000001101111",
    972 => "00111111010010001111100001000011",
    973 => "00111111001010110000010010010111",
    974 => "00111111000111100100110000110111",
    975 => "00111111000111101001010000011101",
    976 => "10111101101001110101110110000010",
    977 => "10111110001101000010011110101110",
    978 => "00111111100011111100100110110001",
    979 => "10111101111001011001001110010101",
    980 => "10111101111001011001001110101001",
    981 => "00111101111001011001001110101001",
    982 => "00111111011111100110001010000000",
    983 => "00111111011111100110001011101111",
    984 => "10111111011111100110001011101111",
    985 => "10111101010000000110010101011000",
    986 => "10111110001001111000000111000100",
    987 => "00111111101001010001001101011000",
    988 => "00111111001010110000010010010111",
    989 => "00111111010001101110000001101111",
    990 => "00111111010010001111100001000011",
    991 => "00111111001010110000010010010111",
    992 => "00111111000111100100110000110111",
    993 => "00111111000111101001010000011101",
    994 => "10111110110000001110110111111010",
    995 => "00111101010111000110010001101001",
    996 => "10111111011011001011101010111100",
    997 => "10111101001110100000110100100110",
    998 => "10111110001001010000000010100000",
    999 => "00111111101001111000110101110011");


  component fsub is
    port (A : in std_logic_vector (31 downto 0);
          B : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          C : out std_logic_vector (31 downto 0));
  end component fsub;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal s_b : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (4 downto 0) of std_logic_vector (31 downto 0);
  signal cc : buff := (others => (others => '0'));
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
  signal i_isRunning : std_logic := 'U';
  signal i_result : std_logic := '1';
begin  -- architecture fsub_tb

  i_fsub : fsub port map (s_a,s_b,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk) is
    variable ss : character;
    variable count : integer := 4;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      case state is
        when "00" =>
          state <= "01";
        when "01" =>
          state <= "11";
        when "11" =>
          state <= "10";
        when others =>
          state <= "00";
      end case;
      s_a <= a_lut (addr);
      s_b <= b_lut (addr);
      cc(conv_integer(state)) <= ans_lut (addr);      
      ccc <= cc (conv_integer (state));
      if i_isRunning = '1' then  -- rising clock edge
        if ccc = c and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 5 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;
  end process ram_loop;

end architecture;
