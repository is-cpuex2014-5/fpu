library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity fsqrt_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity fsqrt_tb;

architecture testbench of fsqrt_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "01000000010100000000000000000000",
    1 => "00111111100000000000000000000001",
    2 => "00111101110011001100110011001101",
    3 => "00111101110100000101100110000111",
    4 => "00111111001010011011001111001110",
    5 => "00111101110110000000111110000011",
    6 => "00111111001000010101010000110100",
    7 => "00111101110101111101101100100101",
    8 => "00111111001000011000001011111000",
    9 => "00111101110101111101110001010101",
    10 => "00111111001000011000000111110000",
    11 => "00111101110101111101110001001110",
    12 => "00111111110001001010010100100100",
    13 => "00111101110011001100110011001101",
    14 => "00111111001011101101000001000010",
    15 => "00111111010110100010111111111100",
    16 => "00111111010101110100101100101100",
    17 => "00111111010101110111110011011100",
    18 => "00111111010101110111100110010010",
    19 => "00111111010101110111100111001100",
    20 => "00111111010101110111100111000110",
    21 => "00111111010101110111100111001100",
    22 => "00111111010101110111100111000110",
    23 => "01000000000111101111000000011000",
    24 => "00111101110011001100110011001101",
    25 => "00111101111011111111000001000101",
    26 => "00111111000101010011011010110100",
    27 => "00111110000110010001011110000011",
    28 => "00111111000110000111101011000010",
    29 => "00111110000110010111111000010110",
    30 => "00111111000110001010001010101100",
    31 => "00111110000110011000001011100110",
    32 => "00111111000110001010010010001100",
    33 => "00111110000110011000001100100000",
    34 => "00111111110001011110100100011100",
    35 => "00111101110011001100110011001101",
    36 => "00111110100010100010100011110001",
    37 => "00111111010010000000000110010000",
    38 => "00111110111011111110010110110110",
    39 => "00111111010110110111001001011010",
    40 => "00111110111100011010001010100000",
    41 => "00111111010110110111111101011100",
    42 => "00111110111100011010001110011000",
    43 => "00111111010110110111111101101100",
    44 => "00111110111100011010001110100101",
    45 => "01000000000010000100011110000010",
    46 => "00111101110011001100110011001101",
    47 => "00111110001000101011000101101010",
    48 => "00111111000111000111101111111000",
    49 => "00111110100000100100111001000101",
    50 => "00111111010000111101110011011100",
    51 => "00111110100001101110011001010010",
    52 => "00111111010001100101110001110110",
    53 => "00111110100001110010000111000011",
    54 => "00111111010001100111101101100010",
    55 => "00111110100001110010010010010110",
    56 => "00111111111010110110110111111010",
    57 => "00111101110011001100110011001101",
    58 => "00111110001000101011000101101100",
    59 => "00111111000111000111101111111010",
    60 => "00111110100000100100111001001001",
    61 => "00111111010000111101110011011100",
    62 => "00111110100001101110011001010011",
    63 => "00111111010001100101110001111110",
    64 => "00111110100001110010000111001001",
    65 => "00111111010001100111101101100100",
    66 => "00111110100001110010010010011001",
    67 => "00111111111010110110110111111101",
    68 => "00111101110011001100110011001101",
    69 => "00111110100010100010100100010100",
    70 => "00111111010010000000000110100100",
    71 => "00111110111011111110010110111101",
    72 => "00111111010110110111001001011010",
    73 => "00111110111100011010001010010110",
    74 => "00111111010110110111111101100010",
    75 => "00111110111100011010001110011101",
    76 => "00111111010110110111111101100010",
    77 => "00111110111100011010001110011101",
    78 => "01000000000010000100011101111111",
    79 => "00111101110011001100110011001101",
    80 => "00111101111011111111000001000110",
    81 => "00111111000101010011011010110101",
    82 => "00111110000110010001011110000100",
    83 => "00111111000110000111101011000011",
    84 => "00111110000110010111111000011000",
    85 => "00111111000110001010001010101110",
    86 => "00111110000110011000001011101000",
    87 => "00111111000110001010010010001110",
    88 => "00111110000110011000001100100010",
    89 => "00111111110001011110100100011110",
    90 => "00111101110011001100110011001101",
    91 => "00111111001011101101100011000110",
    92 => "00111111010110100010111101110110",
    93 => "00111111010101110100101100110000",
    94 => "00111111010101110111110011011000",
    95 => "00111111010101110111100110001110",
    96 => "00111111010101110111100111010100",
    97 => "00111111010101110111100110111100",
    98 => "00111111010101110111100111000110",
    99 => "00111111010101110111100111000100",
    100 => "01000000000111101111000000010111",
    101 => "00111101110011001100110011001101",
    102 => "00111101110100000101100110000111",
    103 => "00111111001010011011001111001110",
    104 => "00111101110110000000111110000011",
    105 => "00111111001000010101010000110100",
    106 => "00111101110101111101101100100101",
    107 => "00111111001000011000001011111000",
    108 => "00111101110101111101110001010101",
    109 => "00111111001000011000000111110000",
    110 => "00111101110101111101110001001110",
    111 => "00111111110001001010010100100100",
    112 => "00111101110011001100110011001101",
    113 => "00111101110100000101100110000110",
    114 => "00111110100010010001000011100000",
    115 => "00111101110100111100001111110001",
    116 => "00111110100010000011010110011001",
    117 => "00111101110100111011101111010000",
    118 => "00111110100010000011011101101111",
    119 => "00111101110100111011101111100010",
    120 => "00111110100010000011011101101100",
    121 => "00111101110100111011101111100010",
    122 => "00111111100101011011000000000000",
    123 => "00111101110011001100110011001101",
    124 => "00111111001011101101000001001000",
    125 => "00111110111011001101000111000001",
    126 => "00111111010110110101100001111000",
    127 => "00111110111100011010000010001101",
    128 => "00111111010110110111111101010110",
    129 => "00111110111100011010001110100101",
    130 => "00111111010110110111111101100110",
    131 => "00111110111100011010001110100010",
    132 => "00111111010110110111111101100100",
    133 => "01000000000010000100011110000000",
    134 => "00111101110011001100110011001101",
    135 => "00111101111011111111000001000101",
    136 => "00111110100001100000100111000111",
    137 => "00111110000001110111010111010001",
    138 => "00111110100010001111111110100000",
    139 => "00111110000001111111101010111100",
    140 => "00111110100010010010011000101010",
    141 => "00111110000010000000000101101100",
    142 => "00111110100010010010100000100011",
    143 => "00111110000010000000000111000100",
    144 => "00111111100110011011000010101110",
    145 => "00111101110011001100110011001101",
    146 => "00111110100010100010100011110001",
    147 => "00111110101111010000110001011100",
    148 => "00111110110100110001011010010000",
    149 => "00111110110110010110001001101001",
    150 => "00111110110110101110110110010010",
    151 => "00111110110110110100101010010011",
    152 => "00111110110110110110000001000011",
    153 => "00111110110110110110010101001101",
    154 => "00111110110110110110011001110101",
    155 => "00111111110101000001100110110011",
    156 => "00111101110011001100110011001101",
    157 => "00111110001000101011000101101010",
    158 => "00111110100100101111101101100110",
    159 => "00111110010101111011100001011110",
    160 => "00111110101010001100011101101001",
    161 => "00111110011000010101100010101110",
    162 => "00111110101011000110100001011111",
    163 => "00111110011000101100100101000111",
    164 => "00111110101011001111000000001011",
    165 => "00111110011000101111111000110100",
    166 => "00111111101011100000011100001000",
    167 => "00111101110011001100110011001101",
    168 => "00111110001000101011000101101100",
    169 => "00111110100100101111101101100111",
    170 => "00111110010101111011100001100111",
    171 => "00111110101010001100011101101000",
    172 => "00111110011000010101100010101111",
    173 => "00111110101011000110100001011111",
    174 => "00111110011000101100100101000111",
    175 => "00111110101011001111000000001011",
    176 => "00111110011000101111111000111000",
    177 => "00111111101011100000011100001010",
    178 => "00111101110011001100110011001101",
    179 => "00111110100010100010100100010100",
    180 => "00111110101111010000110001110101",
    181 => "00111110110100110001011010011001",
    182 => "00111110110110010110001001101001",
    183 => "00111110110110101110110110001101",
    184 => "00111110110110110100101010010000",
    185 => "00111110110110110110000000111001",
    186 => "00111110110110110110010101001011",
    187 => "00111110110110110110011001101100",
    188 => "00111111110101000001100110110000",
    189 => "00111101110011001100110011001101",
    190 => "00111101111011111111000001000110",
    191 => "00111110100001100000100111000111",
    192 => "00111110000001110111010111010010",
    193 => "00111110100010001111111110100000",
    194 => "00111110000001111111101010111101",
    195 => "00111110100010010010011000101010",
    196 => "00111110000010000000000101101100",
    197 => "00111110100010010010100000100011",
    198 => "00111110000010000000000111000101",
    199 => "00111111100110011011000010101110",
    200 => "00111101110011001100110011001101",
    201 => "00111111001011101101100011000110",
    202 => "00111110111011001101001100001000",
    203 => "00111111010110110101100011000110",
    204 => "00111110111100011010000010011100",
    205 => "00111111010110110111111110001100",
    206 => "00111110111100011010001110101010",
    207 => "00111111010110110111111110011010",
    208 => "00111110111100011010001110100101",
    209 => "00111111010110110111111110100100",
    210 => "01000000000010000100011110010010",
    211 => "00111101110011001100110011001101",
    212 => "00111101110100000101100110000111",
    213 => "00111110100010010001000011100000",
    214 => "00111101110100111100001111110010",
    215 => "00111110100010000011010110010111",
    216 => "00111101110100111011101111010001",
    217 => "00111110100010000011011101101100",
    218 => "00111101110100111011101111100010",
    219 => "00111110100010000011011101101100",
    220 => "00111101110100111011101111100010",
    221 => "00111111100101011011000000000000",
    222 => "00111101110011001100110011001101",
    223 => "00111101110100000101100110000111",
    224 => "00111110001000100111000010101011",
    225 => "00111101110100010101111010010001",
    226 => "00111110001000100110001001001001",
    227 => "00111101110100010101111000111100",
    228 => "00111110001000100110001001001110",
    229 => "00111101110100010101111000111100",
    230 => "00111110001000100110001001001110",
    231 => "00111101110100010101111000111100",
    232 => "00111111100001111100100010010100",
    233 => "00111101110011001100110011001101",
    234 => "00111111001011101101000001000010",
    235 => "00111110100001001011000001110011",
    236 => "00111111010001010010111110011000",
    237 => "00111110100001110000010111111101",
    238 => "00111111010001100110110011101100",
    239 => "00111110100001110010001101000110",
    240 => "00111111010001100111110000101010",
    241 => "00111110100001110010010010101010",
    242 => "00111111010001100111110011011110",
    243 => "00111111111010110110111000000100",
    244 => "00111101110011001100110011001101",
    245 => "00111101111011111111000001000101",
    246 => "00111110001000110010000100111000",
    247 => "00111101111110010101110000011000",
    248 => "00111110001001000000000101000000",
    249 => "00111101111110011000110101010100",
    250 => "00111110001001000000011001100000",
    251 => "00111101111110011000111001110101",
    252 => "00111110001001000000011001111101",
    253 => "00111101111110011000111001111010",
    254 => "00111111100010101000000000011110",
    255 => "00111101110011001100110011001101",
    256 => "00111110100010100010100011110001",
    257 => "00111110010100110100110010101000",
    258 => "00111110101001110001000001011110",
    259 => "00111110011000001010011010011110",
    260 => "00111110101011000010011001111110",
    261 => "00111110011000101010111101111100",
    262 => "00111110101011001110011010000110",
    263 => "00111110011000101111101001111000",
    264 => "00111110101011010000001000001010",
    265 => "00111111101011100000011110010000",
    266 => "00111101110011001100110011001101",
    267 => "00111110001000101011000101101010",
    268 => "00111110001011110110000100010100",
    269 => "00111110001100111100110000110000",
    270 => "00111110001101010101011111101010",
    271 => "00111110001101011110001000110011",
    272 => "00111110001101100001001001111111",
    273 => "00111110001101100010001101010110",
    274 => "00111110001101100010100100111100",
    275 => "00111110001101100010101101000110",
    276 => "00111111100100111111000101001111",
    277 => "00111101110011001100110011001101",
    278 => "00111110001000101011000101101100",
    279 => "00111110001011110110000100010100",
    280 => "00111110001100111100110000110011",
    281 => "00111110001101010101011111101100",
    282 => "00111110001101011110001000110110",
    283 => "00111110001101100001001001111110",
    284 => "00111110001101100010001101011010",
    285 => "00111110001101100010100100111110",
    286 => "00111110001101100010101101001100",
    287 => "00111111100100111111000101010000",
    288 => "00111101110011001100110011001101",
    289 => "00111110100010100010100100010100",
    290 => "00111110010100110100110011000000",
    291 => "00111110101001110001000001100100",
    292 => "00111110011000001010011010011100",
    293 => "00111110101011000010011001101110",
    294 => "00111110011000101010111101111010",
    295 => "00111110101011001110011001111101",
    296 => "00111110011000101111101001110110",
    297 => "00111110101011010000000111111110",
    298 => "00111111101011100000011110001100",
    299 => "00111101110011001100110011001101",
    300 => "00111101111011111111000001000110",
    301 => "00111110001000110010000100111000",
    302 => "00111101111110010101110000011001",
    303 => "00111110001001000000000101000000",
    304 => "00111101111110011000110101010100",
    305 => "00111110001001000000011001100000",
    306 => "00111101111110011000111001110110",
    307 => "00111110001001000000011001111101",
    308 => "00111101111110011000111001111100",
    309 => "00111111100010101000000000011110",
    310 => "00111101110011001100110011001101",
    311 => "00111111001011101101100011000110",
    312 => "00111110100001001011000101110100",
    313 => "00111111010001010011000110010110",
    314 => "00111110100001110000011000110000",
    315 => "00111111010001100110111001110110",
    316 => "00111110100001110010001101101100",
    317 => "00111111010001100111110110011110",
    318 => "00111110100001110010010011001101",
    319 => "00111111010001100111111001010110",
    320 => "00111111111010110110111011001001",
    321 => "00111101110011001100110011001101",
    322 => "00111101110100000101100110000111",
    323 => "00111110001000100111000010101011",
    324 => "00111101110100010101111010010001",
    325 => "00111110001000100110001001001001",
    326 => "00111101110100010101111000111100",
    327 => "00111110001000100110001001001110",
    328 => "00111101110100010101111000111100",
    329 => "00111110001000100110001001001110",
    330 => "00111101110100010101111000111100",
    331 => "00111111100001111100100010010100",
    332 => "00111101110011001100110011001101",
    333 => "00111101110100000101100110000110",
    334 => "00111101111011111110110011100100",
    335 => "00111101110100001000001000000010",
    336 => "00111101111011111110110011111001",
    337 => "00111101110100001000001000000010",
    338 => "00111101111011111110110011111001",
    339 => "00111101110100001000001000000010",
    340 => "00111101111011111110110011111001",
    341 => "00111101110100001000001000000010",
    342 => "00111111100000100110110101010110",
    343 => "00111101110011001100110011001101",
    344 => "00111111001011101101000001001000",
    345 => "00111110000110111110011101000001",
    346 => "00111111000110011001100010111101",
    347 => "00111110000110011010000001100100",
    348 => "00111111000110001011000000000010",
    349 => "00111110000110011000010010000011",
    350 => "00111111000110001010010100101110",
    351 => "00111110000110011000001100110110",
    352 => "00111111000110001010010010110001",
    353 => "00111111110001011110100100100100",
    354 => "00111101110011001100110011001101",
    355 => "00111101111011111111000001000101",
    356 => "00111101111100010001111000110101",
    357 => "00111101111100010011001000010010",
    358 => "00111101111100010011001101101001",
    359 => "00111101111100010011001101111101",
    360 => "00111101111100010011001110000000",
    361 => "00111101111100010011001101111110",
    362 => "00111101111100010011001110000000",
    363 => "00111101111100010011001101111110",
    364 => "00111111100001001000110011010110",
    365 => "00111101110011001100110011001101",
    366 => "00111110100010100010100011110001",
    367 => "00111110000010000010111000101000",
    368 => "00111110100010010011010101000100",
    369 => "00111110000010000000010000001101",
    370 => "00111110100010010010100011100111",
    371 => "00111110000010000000000111101001",
    372 => "00111110100010010010100001000100",
    373 => "00111110000010000000000111001100",
    374 => "00111110100010010010100000111011",
    375 => "00111111100110011011000010101110",
    376 => "00111101110011001100110011001101",
    377 => "00111110001000101011000101101010",
    378 => "00111101111110010100001110001111",
    379 => "00111110001000111111111010110011",
    380 => "00111101111110011000110011001000",
    381 => "00111110001001000000011001001111",
    382 => "00111101111110011000111001110101",
    383 => "00111110001001000000011001111010",
    384 => "00111101111110011000111001111110",
    385 => "00111110001001000000011001111100",
    386 => "00111111100010101000000000011110",
    387 => "00111101110011001100110011001101",
    388 => "00111110001000101011000101101100",
    389 => "00111101111110010100001110001111",
    390 => "00111110001000111111111010110100",
    391 => "00111101111110011000110011001000",
    392 => "00111110001001000000011001010001",
    393 => "00111101111110011000111001110110",
    394 => "00111110001001000000011001111101",
    395 => "00111101111110011000111001111110",
    396 => "00111110001001000000011001111100",
    397 => "00111111100010101000000000011110",
    398 => "00111101110011001100110011001101",
    399 => "00111110100010100010100100010100",
    400 => "00111110000010000010111000101111",
    401 => "00111110100010010011010100111110",
    402 => "00111110000010000000010000001100",
    403 => "00111110100010010010100011100001",
    404 => "00111110000010000000000111101000",
    405 => "00111110100010010010100001000010",
    406 => "00111110000010000000000111001011",
    407 => "00111110100010010010100000111000",
    408 => "00111111100110011011000010101110",
    409 => "00111101110011001100110011001101",
    410 => "00111101111011111111000001000110",
    411 => "00111101111100010001111000110101",
    412 => "00111101111100010011001000010011",
    413 => "00111101111100010011001101101001",
    414 => "00111101111100010011001101111111",
    415 => "00111101111100010011001110000000",
    416 => "00111101111100010011001101111111",
    417 => "00111101111100010011001110000000",
    418 => "00111101111100010011001101111111",
    419 => "00111111100001001000110011010110",
    420 => "00111101110011001100110011001101",
    421 => "00111111001011101101100011000110",
    422 => "00111110000110111110100000010101",
    423 => "00111111000110011001101100101000",
    424 => "00111110000110011010000010101110",
    425 => "00111111000110001011001000111001",
    426 => "00111110000110011000010011001000",
    427 => "00111111000110001010011101011000",
    428 => "00111110000110011000001101111000",
    429 => "00111111000110001010011011011010",
    430 => "00111111110001011110101001000000",
    431 => "00111101110011001100110011001101",
    432 => "00111101110100000101100110000111",
    433 => "00111101111011111110110011100100",
    434 => "00111101110100001000001000000010",
    435 => "00111101111011111110110011111001",
    436 => "00111101110100001000001000000010",
    437 => "00111101111011111110110011111001",
    438 => "00111101110100001000001000000010",
    439 => "00111101111011111110110011111001",
    440 => "00111101110100001000001000000010",
    441 => "00111111100000100110110101010110",
    442 => "00111101110011001100110011001101",
    443 => "00111101110100000101100110000111",
    444 => "00111101110100000101101010011010",
    445 => "00111101110100000101101010011010",
    446 => "00111101110100000101101010011010",
    447 => "00111101110100000101101010011010",
    448 => "00111101110100000101101010011010",
    449 => "00111101110100000101101010011010",
    450 => "00111101110100000101101010011010",
    451 => "00111101110100000101101010011010",
    452 => "00111111100000000111000110111010",
    453 => "00111101110011001100110011001101",
    454 => "00111111001011101101000001000010",
    455 => "00111101110110000010110110001110",
    456 => "00111111001000010011100110010010",
    457 => "00111101110101111101101001111000",
    458 => "00111111001000011000001110000000",
    459 => "00111101110101111101110001011001",
    460 => "00111111001000011000000111101110",
    461 => "00111101110101111101110001001111",
    462 => "00111111001000011000000111011110",
    463 => "00111111110001001010010100011010",
    464 => "00111101110011001100110011001101",
    465 => "00111101111011111111000001000101",
    466 => "00111101110100001000001000001001",
    467 => "00111101111011111110110011111000",
    468 => "00111101110100001000001000000010",
    469 => "00111101111011111110110011111000",
    470 => "00111101110100001000001000000010",
    471 => "00111101111011111110110011111000",
    472 => "00111101110100001000001000000010",
    473 => "00111101111011111110110011111000",
    474 => "00111111100000100110110101010110",
    475 => "00111101110011001100110011001101",
    476 => "00111110100010100010100011110001",
    477 => "00111101110100111100111001000011",
    478 => "00111110100010000011001100111111",
    479 => "00111101110100111011101110111011",
    480 => "00111110100010000011011101101100",
    481 => "00111101110100111011101111100010",
    482 => "00111110100010000011011101100111",
    483 => "00111101110100111011101111100010",
    484 => "00111110100010000011011101100111",
    485 => "00111111100101011010111111111110",
    486 => "00111101110011001100110011001101",
    487 => "00111110001000101011000101101010",
    488 => "00111101110100010110000000001110",
    489 => "00111110001000100110001000110010",
    490 => "00111101110100010101111000111100",
    491 => "00111110001000100110001001001100",
    492 => "00111101110100010101111000111100",
    493 => "00111110001000100110001001001100",
    494 => "00111101110100010101111000111100",
    495 => "00111110001000100110001001001100",
    496 => "00111111100001111100100010010100",
    497 => "00111101110011001100110011001101",
    498 => "00111110001000101011000101101100",
    499 => "00111101110100010110000000001110",
    500 => "00111110001000100110001000110110",
    501 => "00111101110100010101111000111100",
    502 => "00111110001000100110001001001110",
    503 => "00111101110100010101111000111100",
    504 => "00111110001000100110001001001110",
    505 => "00111101110100010101111000111100",
    506 => "00111110001000100110001001001110",
    507 => "00111111100001111100100010010100",
    508 => "00111101110011001100110011001101",
    509 => "00111110100010100010100100010100",
    510 => "00111101110100111100111001000100",
    511 => "00111110100010000011001101010111",
    512 => "00111101110100111011101110111100",
    513 => "00111110100010000011011110000011",
    514 => "00111101110100111011101111100100",
    515 => "00111110100010000011011101111100",
    516 => "00111101110100111011101111100011",
    517 => "00111110100010000011011101111100",
    518 => "00111111100101011011000000000100",
    519 => "00111101110011001100110011001101",
    520 => "00111101111011111111000001000110",
    521 => "00111101110100001000001000001001",
    522 => "00111101111011111110110011111001",
    523 => "00111101110100001000001000000010",
    524 => "00111101111011111110110011111001",
    525 => "00111101110100001000001000000010",
    526 => "00111101111011111110110011111001",
    527 => "00111101110100001000001000000010",
    528 => "00111101111011111110110011111001",
    529 => "00111111100000100110110101010110",
    530 => "00111101110011001100110011001101",
    531 => "00111111001011101101100011000110",
    532 => "00111101110110000010110110111111",
    533 => "00111111001000010011111100110100",
    534 => "00111101110101111101101010011101",
    535 => "00111111001000011000100100111010",
    536 => "00111101110101111101110001111110",
    537 => "00111111001000011000011110001010",
    538 => "00111101110101111101110001110011",
    539 => "00111111001000011000011110011110",
    540 => "00111111110001001010011111111100",
    541 => "00111101110011001100110011001101",
    542 => "00111101110100000101100110000111",
    543 => "00111101110100000101101010011010",
    544 => "00111101110100000101101010011010",
    545 => "00111101110100000101101010011010",
    546 => "00111101110100000101101010011010",
    547 => "00111101110100000101101010011010",
    548 => "00111101110100000101101010011010",
    549 => "00111101110100000101101010011010",
    550 => "00111101110100000101101010011010",
    551 => "00111111100000000111000110111010",
    552 => "00111101110011001100110011001101",
    553 => "00111101110100000101100110000110",
    554 => "00111101110100000101101010011001",
    555 => "00111101110100000101101010011010",
    556 => "00111101110100000101101010011010",
    557 => "00111101110100000101101010011010",
    558 => "00111101110100000101101010011010",
    559 => "00111101110100000101101010011010",
    560 => "00111101110100000101101010011010",
    561 => "00111101110100000101101010011010",
    562 => "00111111100000000111000110111010",
    563 => "00111101110011001100110011001101",
    564 => "00111111001011101101000001001000",
    565 => "00111101110110000010110110001100",
    566 => "00111111001000010011100110101000",
    567 => "00111101110101111101101001110111",
    568 => "00111111001000011000001110001000",
    569 => "00111101110101111101110001010111",
    570 => "00111111001000011000000111110100",
    571 => "00111101110101111101110001001101",
    572 => "00111111001000011000000111110000",
    573 => "00111111110001001010010100100100",
    574 => "00111101110011001100110011001101",
    575 => "00111101111011111111000001000101",
    576 => "00111101110100001000001000001000",
    577 => "00111101111011111110110011111000",
    578 => "00111101110100001000001000000010",
    579 => "00111101111011111110110011111000",
    580 => "00111101110100001000001000000010",
    581 => "00111101111011111110110011111000",
    582 => "00111101110100001000001000000010",
    583 => "00111101111011111110110011111000",
    584 => "00111111100000100110110101010110",
    585 => "00111101110011001100110011001101",
    586 => "00111110100010100010100011110001",
    587 => "00111101110100111100111001000010",
    588 => "00111110100010000011001100111111",
    589 => "00111101110100111011101110111010",
    590 => "00111110100010000011011101101100",
    591 => "00111101110100111011101111100010",
    592 => "00111110100010000011011101100111",
    593 => "00111101110100111011101111100010",
    594 => "00111110100010000011011101100111",
    595 => "00111111100101011010111111111110",
    596 => "00111101110011001100110011001101",
    597 => "00111110001000101011000101101010",
    598 => "00111101110100010110000000001101",
    599 => "00111110001000100110001000110010",
    600 => "00111101110100010101111000111011",
    601 => "00111110001000100110001001001100",
    602 => "00111101110100010101111000111100",
    603 => "00111110001000100110001001001100",
    604 => "00111101110100010101111000111100",
    605 => "00111110001000100110001001001100",
    606 => "00111111100001111100100010010100",
    607 => "00111101110011001100110011001101",
    608 => "00111110001000101011000101101100",
    609 => "00111101110100010110000000001101",
    610 => "00111110001000100110001000110110",
    611 => "00111101110100010101111000111011",
    612 => "00111110001000100110001001001110",
    613 => "00111101110100010101111000111100",
    614 => "00111110001000100110001001001110",
    615 => "00111101110100010101111000111100",
    616 => "00111110001000100110001001001110",
    617 => "00111111100001111100100010010100",
    618 => "00111101110011001100110011001101",
    619 => "00111110100010100010100100010100",
    620 => "00111101110100111100111001000011",
    621 => "00111110100010000011001101010111",
    622 => "00111101110100111011101110111010",
    623 => "00111110100010000011011110000011",
    624 => "00111101110100111011101111100010",
    625 => "00111110100010000011011101111111",
    626 => "00111101110100111011101111100010",
    627 => "00111110100010000011011101111111",
    628 => "00111111100101011011000000000100",
    629 => "00111101110011001100110011001101",
    630 => "00111101111011111111000001000110",
    631 => "00111101110100001000001000001000",
    632 => "00111101111011111110110011111010",
    633 => "00111101110100001000001000000010",
    634 => "00111101111011111110110011111001",
    635 => "00111101110100001000001000000010",
    636 => "00111101111011111110110011111001",
    637 => "00111101110100001000001000000010",
    638 => "00111101111011111110110011111001",
    639 => "00111111100000100110110101010110",
    640 => "00111101110011001100110011001101",
    641 => "00111111001011101101100011000110",
    642 => "00111101110110000010110110111101",
    643 => "00111111001000010011111100110100",
    644 => "00111101110101111101101010011011",
    645 => "00111111001000011000100100111010",
    646 => "00111101110101111101110001111100",
    647 => "00111111001000011000011110001000",
    648 => "00111101110101111101110001110001",
    649 => "00111111001000011000011110011110",
    650 => "00111111110001001010011111111100",
    651 => "00111101110011001100110011001101",
    652 => "00111101110100000101100110000111",
    653 => "00111101110100000101101010011001",
    654 => "00111101110100000101101010011010",
    655 => "00111101110100000101101010011010",
    656 => "00111101110100000101101010011010",
    657 => "00111101110100000101101010011010",
    658 => "00111101110100000101101010011010",
    659 => "00111101110100000101101010011010",
    660 => "00111101110100000101101010011010",
    661 => "00111111100000000111000110111010",
    662 => "00111101110011001100110011001101",
    663 => "00111101110100000101100110000111",
    664 => "00111101111011111110110011100010",
    665 => "00111101110100001000001000000010",
    666 => "00111101111011111110110011111000",
    667 => "00111101110100001000001000000010",
    668 => "00111101111011111110110011111000",
    669 => "00111101110100001000001000000010",
    670 => "00111101111011111110110011111000",
    671 => "00111101110100001000001000000010",
    672 => "00111111100000100110110101010110",
    673 => "00111101110011001100110011001101",
    674 => "00111111001011101101000001000010",
    675 => "00111110000110111110011100111110",
    676 => "00111111000110011001100010111110",
    677 => "00111110000110011010000001100010",
    678 => "00111111000110001011000000000010",
    679 => "00111110000110011000010010000000",
    680 => "00111111000110001010010100100010",
    681 => "00111110000110011000001100110010",
    682 => "00111111000110001010010010100100",
    683 => "00111111110001011110100100011101",
    684 => "00111101110011001100110011001101",
    685 => "00111101111011111111000001000101",
    686 => "00111101111100010001111000110011",
    687 => "00111101111100010011001000010010",
    688 => "00111101111100010011001101100111",
    689 => "00111101111100010011001101111100",
    690 => "00111101111100010011001101111110",
    691 => "00111101111100010011001101111110",
    692 => "00111101111100010011001101111110",
    693 => "00111101111100010011001101111110",
    694 => "00111111100001001000110011010110",
    695 => "00111101110011001100110011001101",
    696 => "00111110100010100010100011110001",
    697 => "00111110000010000010111000100110",
    698 => "00111110100010010011010100111111",
    699 => "00111110000010000000010000001011",
    700 => "00111110100010010010100011100100",
    701 => "00111110000010000000000111100111",
    702 => "00111110100010010010100001000011",
    703 => "00111110000010000000000111001010",
    704 => "00111110100010010010100000111010",
    705 => "00111111100110011011000010101110",
    706 => "00111101110011001100110011001101",
    707 => "00111110001000101011000101101010",
    708 => "00111101111110010100001110001101",
    709 => "00111110001000111111111010110011",
    710 => "00111101111110011000110011000100",
    711 => "00111110001001000000011001001111",
    712 => "00111101111110011000111001110010",
    713 => "00111110001001000000011001111001",
    714 => "00111101111110011000111001111011",
    715 => "00111110001001000000011001111011",
    716 => "00111111100010101000000000011101",
    717 => "00111101110011001100110011001101",
    718 => "00111110001000101011000101101100",
    719 => "00111101111110010100001110001110",
    720 => "00111110001000111111111010110100",
    721 => "00111101111110011000110011000101",
    722 => "00111110001001000000011001010001",
    723 => "00111101111110011000111001110010",
    724 => "00111110001001000000011001111100",
    725 => "00111101111110011000111001111010",
    726 => "00111110001001000000011001111110",
    727 => "00111111100010101000000000011110",
    728 => "00111101110011001100110011001101",
    729 => "00111110100010100010100100010100",
    730 => "00111110000010000010111000101100",
    731 => "00111110100010010011010100111111",
    732 => "00111110000010000000010000001011",
    733 => "00111110100010010010100011100000",
    734 => "00111110000010000000000111100110",
    735 => "00111110100010010010100001000010",
    736 => "00111110000010000000000111001001",
    737 => "00111110100010010010100000110111",
    738 => "00111111100110011011000010101101",
    739 => "00111101110011001100110011001101",
    740 => "00111101111011111111000001000110",
    741 => "00111101111100010001111000110011",
    742 => "00111101111100010011001000010100",
    743 => "00111101111100010011001101100110",
    744 => "00111101111100010011001101111110",
    745 => "00111101111100010011001101111110",
    746 => "00111101111100010011001101111111",
    747 => "00111101111100010011001101111110",
    748 => "00111101111100010011001101111111",
    749 => "00111111100001001000110011010110",
    750 => "00111101110011001100110011001101",
    751 => "00111111001011101101100011000110",
    752 => "00111110000110111110100000010010",
    753 => "00111111000110011001101100100110",
    754 => "00111110000110011010000010101011",
    755 => "00111111000110001011001000110110",
    756 => "00111110000110011000010011000101",
    757 => "00111111000110001010011101010110",
    758 => "00111110000110011000001101110101",
    759 => "00111111000110001010011011010110",
    760 => "00111111110001011110101000111110",
    761 => "00111101110011001100110011001101",
    762 => "00111101110100000101100110000111",
    763 => "00111101111011111110110011100010",
    764 => "00111101110100001000001000000010",
    765 => "00111101111011111110110011111000",
    766 => "00111101110100001000001000000010",
    767 => "00111101111011111110110011111000",
    768 => "00111101110100001000001000000010",
    769 => "00111101111011111110110011111000",
    770 => "00111101110100001000001000000010",
    771 => "00111111100000100110110101010110",
    772 => "00111101110011001100110011001101",
    773 => "00111101110100000101100110000110",
    774 => "00111110001000100111000010101000",
    775 => "00111101110100010101111010010000",
    776 => "00111110001000100110001001000111",
    777 => "00111101110100010101111000111100",
    778 => "00111110001000100110001001001100",
    779 => "00111101110100010101111000111100",
    780 => "00111110001000100110001001001100",
    781 => "00111101110100010101111000111100",
    782 => "00111111100001111100100010010100",
    783 => "00111101110011001100110011001101",
    784 => "00111111001011101101000001001000",
    785 => "00111110100001001011000001101111",
    786 => "00111111010001010010111110100010",
    787 => "00111110100001110000010111111110",
    788 => "00111111010001100110110011110010",
    789 => "00111110100001110010001101000101",
    790 => "00111111010001100111110000101000",
    791 => "00111110100001110010010010101000",
    792 => "00111111010001100111110011100100",
    793 => "00111111111010110110111000000110",
    794 => "00111101110011001100110011001101",
    795 => "00111101111011111111000001000101",
    796 => "00111110001000110010000100110100",
    797 => "00111101111110010101110000010111",
    798 => "00111110001001000000000100111110",
    799 => "00111101111110011000110101010011",
    800 => "00111110001001000000011001100000",
    801 => "00111101111110011000111001110101",
    802 => "00111110001001000000011001111010",
    803 => "00111101111110011000111001111011",
    804 => "00111111100010101000000000011101",
    805 => "00111101110011001100110011001101",
    806 => "00111110100010100010100011110001",
    807 => "00111110010100110100110010100110",
    808 => "00111110101001110001000001011101",
    809 => "00111110011000001010011010010110",
    810 => "00111110101011000010011001111001",
    811 => "00111110011000101010111101110110",
    812 => "00111110101011001110011010000111",
    813 => "00111110011000101111101001111000",
    814 => "00111110101011010000001000001010",
    815 => "00111111101011100000011110001111",
    816 => "00111101110011001100110011001101",
    817 => "00111110001000101011000101101010",
    818 => "00111110001011110110000100001111",
    819 => "00111110001100111100110000101110",
    820 => "00111110001101010101011111100110",
    821 => "00111110001101011110001000110010",
    822 => "00111110001101100001001001111100",
    823 => "00111110001101100010001101011000",
    824 => "00111110001101100010100100111011",
    825 => "00111110001101100010101101000110",
    826 => "00111111100100111111000101001110",
    827 => "00111101110011001100110011001101",
    828 => "00111110001000101011000101101100",
    829 => "00111110001011110110000100010000",
    830 => "00111110001100111100110000110000",
    831 => "00111110001101010101011111100111",
    832 => "00111110001101011110001000110100",
    833 => "00111110001101100001001001111110",
    834 => "00111110001101100010001101011010",
    835 => "00111110001101100010100100111001",
    836 => "00111110001101100010101101001010",
    837 => "00111111100100111111000101001111",
    838 => "00111101110011001100110011001101",
    839 => "00111110100010100010100100010100",
    840 => "00111110010100110100110010111011",
    841 => "00111110101001110001000001100001",
    842 => "00111110011000001010011010011010",
    843 => "00111110101011000010011001101100",
    844 => "00111110011000101010111101110110",
    845 => "00111110101011001110011001111011",
    846 => "00111110011000101111101001110010",
    847 => "00111110101011010000000111111001",
    848 => "00111111101011100000011110001010",
    849 => "00111101110011001100110011001101",
    850 => "00111101111011111111000001000110",
    851 => "00111110001000110010000100110100",
    852 => "00111101111110010101110000011000",
    853 => "00111110001001000000000100111110",
    854 => "00111101111110011000110101010100",
    855 => "00111110001001000000011001100000",
    856 => "00111101111110011000111001110110",
    857 => "00111110001001000000011001111010",
    858 => "00111101111110011000111001111100",
    859 => "00111111100010101000000000011110",
    860 => "00111101110011001100110011001101",
    861 => "00111111001011101101100011000110",
    862 => "00111110100001001011000101110010",
    863 => "00111111010001010011000110010100",
    864 => "00111110100001110000011000101011",
    865 => "00111111010001100110111001110010",
    866 => "00111110100001110010001101101000",
    867 => "00111111010001100111110110011000",
    868 => "00111110100001110010010011001010",
    869 => "00111111010001100111111001010000",
    870 => "00111111111010110110111011000110",
    871 => "00111101110011001100110011001101",
    872 => "00111101110100000101100110000111",
    873 => "00111110001000100111000010101000",
    874 => "00111101110100010101111010010001",
    875 => "00111110001000100110001001000111",
    876 => "00111101110100010101111000111100",
    877 => "00111110001000100110001001001100",
    878 => "00111101110100010101111000111100",
    879 => "00111110001000100110001001001100",
    880 => "00111101110100010101111000111100",
    881 => "00111111100001111100100010010100",
    882 => "00111101110011001100110011001101",
    883 => "00111101110100000101100110000111",
    884 => "00111110100010010001000011111001",
    885 => "00111101110100111100001111110010",
    886 => "00111110100010000011010110101000",
    887 => "00111101110100111011101111010010",
    888 => "00111110100010000011011101111111",
    889 => "00111101110100111011101111100011",
    890 => "00111110100010000011011101111100",
    891 => "00111101110100111011101111100011",
    892 => "00111111100101011011000000000100",
    893 => "00111101110011001100110011001101",
    894 => "00111111001011101101000001000010",
    895 => "00111110111011001101000110111001",
    896 => "00111111010110110101100001110010",
    897 => "00111110111100011010000010000001",
    898 => "00111111010110110111111101000100",
    899 => "00111110111100011010001110011011",
    900 => "00111111010110110111111101011010",
    901 => "00111110111100011010001110011000",
    902 => "00111111010110110111111101100100",
    903 => "01000000000010000100011110000000",
    904 => "00111101110011001100110011001101",
    905 => "00111101111011111111000001000101",
    906 => "00111110100001100000100111000111",
    907 => "00111110000001110111010111010001",
    908 => "00111110100010001111111110011001",
    909 => "00111110000001111111101010111100",
    910 => "00111110100010010010011000100110",
    911 => "00111110000010000000000101101100",
    912 => "00111110100010010010100000011101",
    913 => "00111110000010000000000111000011",
    914 => "00111111100110011011000010101100",
    915 => "00111101110011001100110011001101",
    916 => "00111110100010100010100011110001",
    917 => "00111110101111010000110001010110",
    918 => "00111110110100110001011010001100",
    919 => "00111110110110010110001001100000",
    920 => "00111110110110101110110110010010",
    921 => "00111110110110110100101010001110",
    922 => "00111110110110110110000001000000",
    923 => "00111110110110110110010100111101",
    924 => "00111110110110110110011001110000",
    925 => "00111111110101000001100110101110",
    926 => "00111101110011001100110011001101",
    927 => "00111110001000101011000101101010",
    928 => "00111110100100101111101101011101",
    929 => "00111110010101111011100001011010",
    930 => "00111110101010001100011101011101",
    931 => "00111110011000010101100010100110",
    932 => "00111110101011000110100001000110",
    933 => "00111110011000101100100100111000",
    934 => "00111110101011001110111111110000",
    935 => "00111110011000101111111000100100",
    936 => "00111111101011100000011100000000",
    937 => "00111101110011001100110011001101",
    938 => "00111110001000101011000101101100",
    939 => "00111110100100101111101101011110",
    940 => "00111110010101111011100001100000",
    941 => "00111110101010001100011101011100",
    942 => "00111110011000010101100010101100",
    943 => "00111110101011000110100001001011",
    944 => "00111110011000101100100100111111",
    945 => "00111110101011001110111111110100",
    946 => "00111110011000101111111000101010",
    947 => "00111111101011100000011100000010",
    948 => "00111101110011001100110011001101",
    949 => "00111110100010100010100100010100",
    950 => "00111110101111010000110001101111",
    951 => "00111110110100110001011010010111",
    952 => "00111110110110010110001001011011",
    953 => "00111110110110101110110110001101",
    954 => "00111110110110110100101010001001",
    955 => "00111110110110110110000000111001",
    956 => "00111110110110110110010100111111",
    957 => "00111110110110110110011001101010",
    958 => "00111111110101000001100110101110",
    959 => "00111101110011001100110011001101",
    960 => "00111101111011111111000001000110",
    961 => "00111110100001100000100111001000",
    962 => "00111110000001110111010111010011",
    963 => "00111110100010001111111110011010",
    964 => "00111110000001111111101010111100",
    965 => "00111110100010010010011000100110",
    966 => "00111110000010000000000101101100",
    967 => "00111110100010010010100000011101",
    968 => "00111110000010000000000111000101",
    969 => "00111111100110011011000010101101",
    970 => "00111101110011001100110011001101",
    971 => "00111111001011101101100011000110",
    972 => "00111110111011001101001011111010",
    973 => "00111111010110110101100011000110",
    974 => "00111110111100011010000010001101",
    975 => "00111111010110110111111110001010",
    976 => "00111110111100011010001110011101",
    977 => "00111111010110110111111110011100",
    978 => "00111110111100011010001110011101",
    979 => "00111111010110110111111110011100",
    980 => "01000000000010000100011110001110",
    981 => "00111101110011001100110011001101",
    982 => "00111101110100000101100110000111",
    983 => "00111110100010010001000011111001",
    984 => "00111101110100111100001111110010",
    985 => "00111110100010000011010110101000",
    986 => "00111101110100111011101111010010",
    987 => "00111110100010000011011101111111",
    988 => "00111101110100111011101111100011",
    989 => "00111110100010000011011101111100",
    990 => "00111101110100111011101111100011",
    991 => "00111111100101011011000000000100",
    992 => "00111101110011001100110011001101",
    993 => "00111101110100000101100110000110",
    994 => "00111111001010011011101100111010",
    995 => "00111101110110000000111110101110",
    996 => "00111111001000010101100111001100",
    997 => "00111101110101111101101101001000",
    998 => "00111111001000011000100010101000",
    999 => "00111101110101111101110001111000");

  constant ans_lut : lut := (
    0 => "00111111111001101100000101011010",
    1 => "00111111100000000000000000000000",
    2 => "00111110101000011110100010011011",
    3 => "00111110101000110100111001000100",
    4 => "00111111010100000110111010001000",
    5 => "00111110101001100100110011011001",
    6 => "00111111010010110011100101111001",
    7 => "00111110101001100011100010110001",
    8 => "00111111010010110101011011101100",
    9 => "00111110101001100011100100100110",
    10 => "00111111010010110101011001000110",
    11 => "00111110101001100011100100100011",
    12 => "00111111100111101010011100000000",
    13 => "00111110101000011110100010011011",
    14 => "00111111010100111000110000011011",
    15 => "00111111011011000101011010110101",
    16 => "00111111011010101100010000100110",
    17 => "00111111011010101101111100111100",
    18 => "00111111011010101101110101110001",
    19 => "00111111011010101101110110010000",
    20 => "00111111011010101101110110001101",
    21 => "00111111011010101101110110010000",
    22 => "00111111011010101101110110001101",
    23 => "00111111110010011011011010000000",
    24 => "00111110101000011110100010011011",
    25 => "00111110101011110011111110101111",
    26 => "00111111010000110111000111100100",
    27 => "00111110110001011111011111101100",
    28 => "00111111010001011001001001111001",
    29 => "00111110110001100011101000110101",
    30 => "00111111010001011010110001010011",
    31 => "00111110110001100011110101010000",
    32 => "00111111010001011010110110001010",
    33 => "00111110110001100011110101110101",
    34 => "00111111100111110010100101111011",
    35 => "00111110101000011110100010011011",
    36 => "00111111000001001111101110100011",
    37 => "00111111011000100100011100010010",
    38 => "00111111001011110011101111010100",
    39 => "00111111011011010000010100001101",
    40 => "00111111001011111101111000001000",
    41 => "00111111011011010000110000010011",
    42 => "00111111001011111101111001100010",
    43 => "00111111011011010000110000011100",
    44 => "00111111001011111101111001100111",
    45 => "00111111101110101100100000101111",
    46 => "00111110101000011110100010011011",
    47 => "00111110110011000001010011110110",
    48 => "00111111010010000010011001011110",
    49 => "00111111000000010010010111010001",
    50 => "00111111010111111110101111101010",
    51 => "00111111000000110110011110010001",
    52 => "00111111011000010101100001011111",
    53 => "00111111000000111000010010000001",
    54 => "00111111011000010110100111101111",
    55 => "00111111000000111000010111100001",
    56 => "00111111101011011001100000100101",
    57 => "00111110101000011110100010011011",
    58 => "00111110110011000001010011110111",
    59 => "00111111010010000010011001011111",
    60 => "00111111000000010010010111010011",
    61 => "00111111010111111110101111101010",
    62 => "00111111000000110110011110010010",
    63 => "00111111011000010101100001100011",
    64 => "00111111000000111000010010000100",
    65 => "00111111011000010110100111110000",
    66 => "00111111000000111000010111100011",
    67 => "00111111101011011001100000100110",
    68 => "00111110101000011110100010011011",
    69 => "00111111000001001111101110110100",
    70 => "00111111011000100100011100011101",
    71 => "00111111001011110011101111010111",
    72 => "00111111011011010000010100001101",
    73 => "00111111001011111101111000000100",
    74 => "00111111011011010000110000010110",
    75 => "00111111001011111101111001100100",
    76 => "00111111011011010000110000010110",
    77 => "00111111001011111101111001100100",
    78 => "00111111101110101100100000101101",
    79 => "00111110101000011110100010011011",
    80 => "00111110101011110011111110110000",
    81 => "00111111010000110111000111100101",
    82 => "00111110110001011111011111101101",
    83 => "00111111010001011001001001111010",
    84 => "00111110110001100011101000110110",
    85 => "00111111010001011010110001010100",
    86 => "00111110110001100011110101010001",
    87 => "00111111010001011010110110001011",
    88 => "00111110110001100011110101110111",
    89 => "00111111100111110010100101111011",
    90 => "00111110101000011110100010011011",
    91 => "00111111010100111001000101000010",
    92 => "00111111011011000101011001101100",
    93 => "00111111011010101100010000101000",
    94 => "00111111011010101101111100111010",
    95 => "00111111011010101101110101101111",
    96 => "00111111011010101101110110010101",
    97 => "00111111011010101101110110001000",
    98 => "00111111011010101101110110001101",
    99 => "00111111011010101101110110001100",
    100 => "00111111110010011011011001111111",
    101 => "00111110101000011110100010011011",
    102 => "00111110101000110100111001000100",
    103 => "00111111010100000110111010001000",
    104 => "00111110101001100100110011011001",
    105 => "00111111010010110011100101111001",
    106 => "00111110101001100011100010110001",
    107 => "00111111010010110101011011101100",
    108 => "00111110101001100011100100100110",
    109 => "00111111010010110101011001000110",
    110 => "00111110101001100011100100100011",
    111 => "00111111100111101010011100000000",
    112 => "00111110101000011110100010011011",
    113 => "00111110101000110100111001000100",
    114 => "00111111000001000111010010010110",
    115 => "00111110101001001010001110001111",
    116 => "00111111000001000000101001111000",
    117 => "00111110101001001010000001100110",
    118 => "00111111000001000000101101011100",
    119 => "00111110101001001010000001101101",
    120 => "00111111000001000000101101011010",
    121 => "00111110101001001010000001101101",
    122 => "00111111100010100110101101101110",
    123 => "00111110101000011110100010011011",
    124 => "00111111010100111000110000011111",
    125 => "00111111001011100001101100011110",
    126 => "00111111011011001111011100010010",
    127 => "00111111001011111101110101000111",
    128 => "00111111011011010000110000010000",
    129 => "00111111001011111101111001100111",
    130 => "00111111011011010000110000011001",
    131 => "00111111001011111101111001100110",
    132 => "00111111011011010000110000011000",
    133 => "00111111101110101100100000101110",
    134 => "00111110101000011110100010011011",
    135 => "00111110101011110011111110101111",
    136 => "00111111000000101111101111111011",
    137 => "00111110101110100011100001000101",
    138 => "00111111000001000110110001000000",
    139 => "00111110101110101001001110001100",
    140 => "00111111000001000111111011011110",
    141 => "00111110101110101001100000100010",
    142 => "00111111000001000111111111010010",
    143 => "00111110101110101001100001011111",
    144 => "00111111100011000100001000010100",
    145 => "00111110101000011110100010011011",
    146 => "00111111000001001111101110100011",
    147 => "00111111000110111000111011000001",
    148 => "00111111001001000110000000011011",
    149 => "00111111001001101100111100010011",
    150 => "00111111001001110110011001101011",
    151 => "00111111001001111000100111110101",
    152 => "00111111001001111001001000111110",
    153 => "00111111001001111001010000101011",
    154 => "00111111001001111001010010011100",
    155 => "00111111101001001100010011100010",
    156 => "00111110101000011110100010011011",
    157 => "00111110110011000001010011110110",
    158 => "00111111000010010010100110111100",
    159 => "00111110111010101111111110101000",
    160 => "00111111000100101111101101100100",
    161 => "00111110111100000010111101000111",
    162 => "00111111000101001000110110111011",
    163 => "00111110111100001111001101100110",
    164 => "00111111000101001100100000100011",
    165 => "00111110111100010000111110000010",
    166 => "00111111100101010011111111110101",
    167 => "00111110101000011110100010011011",
    168 => "00111110110011000001010011110111",
    169 => "00111111000010010010100110111101",
    170 => "00111110111010101111111110101101",
    171 => "00111111000100101111101101100011",
    172 => "00111110111100000010111101000111",
    173 => "00111111000101001000110110111011",
    174 => "00111110111100001111001101100110",
    175 => "00111111000101001100100000100011",
    176 => "00111110111100010000111110000100",
    177 => "00111111100101010011111111110110",
    178 => "00111110101000011110100010011011",
    179 => "00111111000001001111101110110100",
    180 => "00111111000110111000111011001011",
    181 => "00111111001001000110000000011111",
    182 => "00111111001001101100111100010011",
    183 => "00111111001001110110011001101001",
    184 => "00111111001001111000100111110100",
    185 => "00111111001001111001001000111010",
    186 => "00111111001001111001010000101010",
    187 => "00111111001001111001010010011000",
    188 => "00111111101001001100010011100001",
    189 => "00111110101000011110100010011011",
    190 => "00111110101011110011111110110000",
    191 => "00111111000000101111101111111011",
    192 => "00111110101110100011100001000101",
    193 => "00111111000001000110110001000000",
    194 => "00111110101110101001001110001100",
    195 => "00111111000001000111111011011110",
    196 => "00111110101110101001100000100010",
    197 => "00111111000001000111111111010010",
    198 => "00111110101110101001100001011111",
    199 => "00111111100011000100001000010100",
    200 => "00111110101000011110100010011011",
    201 => "00111111010100111001000101000010",
    202 => "00111111001011100001101110010110",
    203 => "00111111011011001111011100111100",
    204 => "00111111001011111101110101001100",
    205 => "00111111011011010000110000101101",
    206 => "00111111001011111101111001101001",
    207 => "00111111011011010000110000110101",
    208 => "00111111001011111101111001100111",
    209 => "00111111011011010000110000111010",
    210 => "00111111101110101100100000111010",
    211 => "00111110101000011110100010011011",
    212 => "00111110101000110100111001000100",
    213 => "00111111000001000111010010010110",
    214 => "00111110101001001010001110010000",
    215 => "00111111000001000000101001110111",
    216 => "00111110101001001010000001100111",
    217 => "00111111000001000000101101011010",
    218 => "00111110101001001010000001101101",
    219 => "00111111000001000000101101011010",
    220 => "00111110101001001010000001101101",
    221 => "00111111100010100110101101101110",
    222 => "00111110101000011110100010011011",
    223 => "00111110101000110100111001000100",
    224 => "00111110110010111110110001010110",
    225 => "00111110101000111011010001110001",
    226 => "00111110110010111110001101001110",
    227 => "00111110101000111011010001010000",
    228 => "00111110110010111110001101010001",
    229 => "00111110101000111011010001010000",
    230 => "00111110110010111110001101010001",
    231 => "00111110101000111011010001010000",
    232 => "00111111100000111101010110010110",
    233 => "00111110101000011110100010011011",
    234 => "00111111010100111000110000011011",
    235 => "00111111000000100101001011010011",
    236 => "00111111011000001010110100111000",
    237 => "00111111000000110111011011111101",
    238 => "00111111011000010110000110111000",
    239 => "00111111000000111000010100111110",
    240 => "00111111011000010110101001100001",
    241 => "00111111000000111000010111101011",
    242 => "00111111011000010110101011000111",
    243 => "00111111101011011001100000101000",
    244 => "00111110101000011110100010011011",
    245 => "00111110101011110011111110101111",
    246 => "00111110110011000101101100001001",
    247 => "00111110101100101010011111111110",
    248 => "00111110110011001110011100101101",
    249 => "00111110101100101011100110100000",
    250 => "00111110110011001110101001100000",
    251 => "00111110101100101011101000001000",
    252 => "00111110110011001110101001110010",
    253 => "00111110101100101011101000001001",
    254 => "00111111100001010010010110010010",
    255 => "00111110101000011110100010011011",
    256 => "00111111000001001111101110100011",
    257 => "00111110111010001001010000001010",
    258 => "00111111000100100011101110111011",
    259 => "00111110111011111101000001001111",
    260 => "00111111000101000111000101010111",
    261 => "00111110111100001110010110110001",
    262 => "00111111000101001100010000001010",
    263 => "00111110111100010000110110000110",
    264 => "00111111000101001100111111100001",
    265 => "00111111100101010100000000110000",
    266 => "00111110101000011110100010011011",
    267 => "00111110110011000001010011110110",
    268 => "00111110110100111110001110101001",
    269 => "00111110110101101000101010110100",
    270 => "00111110110101110111011001001011",
    271 => "00111110110101111100100001100010",
    272 => "00111110110101111110010100000111",
    273 => "00111110110101111110111100000010",
    274 => "00111110110101111111001010000010",
    275 => "00111110110101111111001110110111",
    276 => "00111111100010011001110001001011",
    277 => "00111110101000011110100010011011",
    278 => "00111110110011000001010011110111",
    279 => "00111110110100111110001110101001",
    280 => "00111110110101101000101010110110",
    281 => "00111110110101110111011001001100",
    282 => "00111110110101111100100001100100",
    283 => "00111110110101111110010100000110",
    284 => "00111110110101111110111100000101",
    285 => "00111110110101111111001010000011",
    286 => "00111110110101111111001110111011",
    287 => "00111111100010011001110001001011",
    288 => "00111110101000011110100010011011",
    289 => "00111111000001001111101110110100",
    290 => "00111110111010001001010000010111",
    291 => "00111111000100100011101110111101",
    292 => "00111110111011111101000001001110",
    293 => "00111111000101000111000101010000",
    294 => "00111110111100001110010110110000",
    295 => "00111111000101001100010000000110",
    296 => "00111110111100010000110110000101",
    297 => "00111111000101001100111111011100",
    298 => "00111111100101010100000000101110",
    299 => "00111110101000011110100010011011",
    300 => "00111110101011110011111110110000",
    301 => "00111110110011000101101100001001",
    302 => "00111110101100101010011111111110",
    303 => "00111110110011001110011100101101",
    304 => "00111110101100101011100110100000",
    305 => "00111110110011001110101001100000",
    306 => "00111110101100101011101000001000",
    307 => "00111110110011001110101001110010",
    308 => "00111110101100101011101000001010",
    309 => "00111111100001010010010110010010",
    310 => "00111110101000011110100010011011",
    311 => "00111111010100111001000101000010",
    312 => "00111111000000100101001101010001",
    313 => "00111111011000001010111001011011",
    314 => "00111111000000110111011100010110",
    315 => "00111111011000010110001010011000",
    316 => "00111111000000111000010101010000",
    317 => "00111111011000010110101100110100",
    318 => "00111111000000111000010111111100",
    319 => "00111111011000010110101110011101",
    320 => "00111111101011011001100001110001",
    321 => "00111110101000011110100010011011",
    322 => "00111110101000110100111001000100",
    323 => "00111110110010111110110001010110",
    324 => "00111110101000111011010001110001",
    325 => "00111110110010111110001101001110",
    326 => "00111110101000111011010001010000",
    327 => "00111110110010111110001101010001",
    328 => "00111110101000111011010001010000",
    329 => "00111110110010111110001101010001",
    330 => "00111110101000111011010001010000",
    331 => "00111111100000111101010110010110",
    332 => "00111110101000011110100010011011",
    333 => "00111110101000110100111001000100",
    334 => "00111110101011110011111001110011",
    335 => "00111110101000110101111000100001",
    336 => "00111110101011110011111001111011",
    337 => "00111110101000110101111000100001",
    338 => "00111110101011110011111001111011",
    339 => "00111110101000110101111000100001",
    340 => "00111110101011110011111001111011",
    341 => "00111110101000110101111000100001",
    342 => "00111111100000010011010100110101",
    343 => "00111110101000011110100010011011",
    344 => "00111111010100111000110000011111",
    345 => "00111110110001111100011100101011",
    346 => "00111111010001100100101101101000",
    347 => "00111110110001100101000001011001",
    348 => "00111111010001011011010011110110",
    349 => "00111110110001100011111001011010",
    350 => "00111111010001011010110111110011",
    351 => "00111110110001100011110110000100",
    352 => "00111111010001011010110110100010",
    353 => "00111111100111110010100101111110",
    354 => "00111110101000011110100010011011",
    355 => "00111110101011110011111110101111",
    356 => "00111110101011111010110111010001",
    357 => "00111110101011111011010100001101",
    358 => "00111110101011111011010110001010",
    359 => "00111110101011111011010110010001",
    360 => "00111110101011111011010110010010",
    361 => "00111110101011111011010110010010",
    362 => "00111110101011111011010110010010",
    363 => "00111110101011111011010110010010",
    364 => "00111111100000100100000101010100",
    365 => "00111110101000011110100010011011",
    366 => "00111111000001001111101110100011",
    367 => "00111110101110101011011011001111",
    368 => "00111111000001001000011000101010",
    369 => "00111110101110101001100111110000",
    370 => "00111111000001001000000000110001",
    371 => "00111110101110101001100001111000",
    372 => "00111111000001000111111111100010",
    373 => "00111110101110101001100001100100",
    374 => "00111111000001000111111111011110",
    375 => "00111111100011000100001000010100",
    376 => "00111110101000011110100010011011",
    377 => "00111110110011000001010011110110",
    378 => "00111110101100101001111100110100",
    379 => "00111110110011001110010110010101",
    380 => "00111110101100101011100101101110",
    381 => "00111110110011001110101001010110",
    382 => "00111110101100101011101000001000",
    383 => "00111110110011001110101001110000",
    384 => "00111110101100101011101000001011",
    385 => "00111110110011001110101001110010",
    386 => "00111111100001010010010110010010",
    387 => "00111110101000011110100010011011",
    388 => "00111110110011000001010011110111",
    389 => "00111110101100101001111100110100",
    390 => "00111110110011001110010110010110",
    391 => "00111110101100101011100101101110",
    392 => "00111110110011001110101001010111",
    393 => "00111110101100101011101000001000",
    394 => "00111110110011001110101001110010",
    395 => "00111110101100101011101000001011",
    396 => "00111110110011001110101001110010",
    397 => "00111111100001010010010110010010",
    398 => "00111110101000011110100010011011",
    399 => "00111111000001001111101110110100",
    400 => "00111110101110101011011011010100",
    401 => "00111111000001001000011000100111",
    402 => "00111110101110101001100111101111",
    403 => "00111111000001001000000000101110",
    404 => "00111110101110101001100001110111",
    405 => "00111111000001000111111111100001",
    406 => "00111110101110101001100001100011",
    407 => "00111111000001000111111111011101",
    408 => "00111111100011000100001000010100",
    409 => "00111110101000011110100010011011",
    410 => "00111110101011110011111110110000",
    411 => "00111110101011111010110111010001",
    412 => "00111110101011111011010100001101",
    413 => "00111110101011111011010110001010",
    414 => "00111110101011111011010110010010",
    415 => "00111110101011111011010110010010",
    416 => "00111110101011111011010110010010",
    417 => "00111110101011111011010110010010",
    418 => "00111110101011111011010110010010",
    419 => "00111111100000100100000101010100",
    420 => "00111110101000011110100010011011",
    421 => "00111111010100111001000101000010",
    422 => "00111110110001111100011110110011",
    423 => "00111111010001100100110011111000",
    424 => "00111110110001100101000010001001",
    425 => "00111111010001011011011001100101",
    426 => "00111110110001100011111010000111",
    427 => "00111111010001011010111101011001",
    428 => "00111110110001100011110110101110",
    429 => "00111111010001011010111100001000",
    430 => "00111111100111110010100111110000",
    431 => "00111110101000011110100010011011",
    432 => "00111110101000110100111001000100",
    433 => "00111110101011110011111001110011",
    434 => "00111110101000110101111000100001",
    435 => "00111110101011110011111001111011",
    436 => "00111110101000110101111000100001",
    437 => "00111110101011110011111001111011",
    438 => "00111110101000110101111000100001",
    439 => "00111110101011110011111001111011",
    440 => "00111110101000110101111000100001",
    441 => "00111111100000010011010100110101",
    442 => "00111110101000011110100010011011",
    443 => "00111110101000110100111001000100",
    444 => "00111110101000110100111010110000",
    445 => "00111110101000110100111010110000",
    446 => "00111110101000110100111010110000",
    447 => "00111110101000110100111010110000",
    448 => "00111110101000110100111010110000",
    449 => "00111110101000110100111010110000",
    450 => "00111110101000110100111010110000",
    451 => "00111110101000110100111010110000",
    452 => "00111111100000000011100011010000",
    453 => "00111110101000011110100010011011",
    454 => "00111111010100111000110000011011",
    455 => "00111110101001100101100001101001",
    456 => "00111111010010110010100010110011",
    457 => "00111110101001100011100001101110",
    458 => "00111111010010110101011101000010",
    459 => "00111110101001100011100100100111",
    460 => "00111111010010110101011001000101",
    461 => "00111110101001100011100100100100",
    462 => "00111111010010110101011000111011",
    463 => "00111111100111101010011011111100",
    464 => "00111110101000011110100010011011",
    465 => "00111110101011110011111110101111",
    466 => "00111110101000110101111000100100",
    467 => "00111110101011110011111001111011",
    468 => "00111110101000110101111000100001",
    469 => "00111110101011110011111001111011",
    470 => "00111110101000110101111000100001",
    471 => "00111110101011110011111001111011",
    472 => "00111110101000110101111000100001",
    473 => "00111110101011110011111001111011",
    474 => "00111111100000010011010100110101",
    475 => "00111110101000011110100010011011",
    476 => "00111111000001001111101110100011",
    477 => "00111110101001001010011110010010",
    478 => "00111111000001000000100101010100",
    479 => "00111110101001001010000001011110",
    480 => "00111111000001000000101101011010",
    481 => "00111110101001001010000001101101",
    482 => "00111111000001000000101101011000",
    483 => "00111110101001001010000001101101",
    484 => "00111111000001000000101101011000",
    485 => "00111111100010100110101101101101",
    486 => "00111110101000011110100010011011",
    487 => "00111110110011000001010011110110",
    488 => "00111110101000111011010100000110",
    489 => "00111110110010111110001101000000",
    490 => "00111110101000111011010001010000",
    491 => "00111110110010111110001101010000",
    492 => "00111110101000111011010001010000",
    493 => "00111110110010111110001101010000",
    494 => "00111110101000111011010001010000",
    495 => "00111110110010111110001101010000",
    496 => "00111111100000111101010110010110",
    497 => "00111110101000011110100010011011",
    498 => "00111110110011000001010011110111",
    499 => "00111110101000111011010100000110",
    500 => "00111110110010111110001101000010",
    501 => "00111110101000111011010001010000",
    502 => "00111110110010111110001101010001",
    503 => "00111110101000111011010001010000",
    504 => "00111110110010111110001101010001",
    505 => "00111110101000111011010001010000",
    506 => "00111110110010111110001101010001",
    507 => "00111111100000111101010110010110",
    508 => "00111110101000011110100010011011",
    509 => "00111111000001001111101110110100",
    510 => "00111110101001001010011110010010",
    511 => "00111111000001000000100101100000",
    512 => "00111110101001001010000001011110",
    513 => "00111111000001000000101101100101",
    514 => "00111110101001001010000001101110",
    515 => "00111111000001000000101101100010",
    516 => "00111110101001001010000001101110",
    517 => "00111111000001000000101101100010",
    518 => "00111111100010100110101101110000",
    519 => "00111110101000011110100010011011",
    520 => "00111110101011110011111110110000",
    521 => "00111110101000110101111000100100",
    522 => "00111110101011110011111001111011",
    523 => "00111110101000110101111000100001",
    524 => "00111110101011110011111001111011",
    525 => "00111110101000110101111000100001",
    526 => "00111110101011110011111001111011",
    527 => "00111110101000110101111000100001",
    528 => "00111110101011110011111001111011",
    529 => "00111111100000010011010100110101",
    530 => "00111110101000011110100010011011",
    531 => "00111111010100111001000101000010",
    532 => "00111110101001100101100001111011",
    533 => "00111111010010110010110001000000",
    534 => "00111110101001100011100001111100",
    535 => "00111111010010110101101011011100",
    536 => "00111110101001100011100100110110",
    537 => "00111111010010110101100111001100",
    538 => "00111110101001100011100100110001",
    539 => "00111111010010110101100111011001",
    540 => "00111111100111101010100000100110",
    541 => "00111110101000011110100010011011",
    542 => "00111110101000110100111001000100",
    543 => "00111110101000110100111010110000",
    544 => "00111110101000110100111010110000",
    545 => "00111110101000110100111010110000",
    546 => "00111110101000110100111010110000",
    547 => "00111110101000110100111010110000",
    548 => "00111110101000110100111010110000",
    549 => "00111110101000110100111010110000",
    550 => "00111110101000110100111010110000",
    551 => "00111111100000000011100011010000",
    552 => "00111110101000011110100010011011",
    553 => "00111110101000110100111001000100",
    554 => "00111110101000110100111010110000",
    555 => "00111110101000110100111010110000",
    556 => "00111110101000110100111010110000",
    557 => "00111110101000110100111010110000",
    558 => "00111110101000110100111010110000",
    559 => "00111110101000110100111010110000",
    560 => "00111110101000110100111010110000",
    561 => "00111110101000110100111010110000",
    562 => "00111111100000000011100011010000",
    563 => "00111110101000011110100010011011",
    564 => "00111111010100111000110000011111",
    565 => "00111110101001100101100001101000",
    566 => "00111111010010110010100011000001",
    567 => "00111110101001100011100001101110",
    568 => "00111111010010110101011101000111",
    569 => "00111110101001100011100100100111",
    570 => "00111111010010110101011001001001",
    571 => "00111110101001100011100100100011",
    572 => "00111111010010110101011001000110",
    573 => "00111111100111101010011100000000",
    574 => "00111110101000011110100010011011",
    575 => "00111110101011110011111110101111",
    576 => "00111110101000110101111000100011",
    577 => "00111110101011110011111001111011",
    578 => "00111110101000110101111000100001",
    579 => "00111110101011110011111001111011",
    580 => "00111110101000110101111000100001",
    581 => "00111110101011110011111001111011",
    582 => "00111110101000110101111000100001",
    583 => "00111110101011110011111001111011",
    584 => "00111111100000010011010100110101",
    585 => "00111110101000011110100010011011",
    586 => "00111111000001001111101110100011",
    587 => "00111110101001001010011110010010",
    588 => "00111111000001000000100101010100",
    589 => "00111110101001001010000001011110",
    590 => "00111111000001000000101101011010",
    591 => "00111110101001001010000001101101",
    592 => "00111111000001000000101101011000",
    593 => "00111110101001001010000001101101",
    594 => "00111111000001000000101101011000",
    595 => "00111111100010100110101101101101",
    596 => "00111110101000011110100010011011",
    597 => "00111110110011000001010011110110",
    598 => "00111110101000111011010100000110",
    599 => "00111110110010111110001101000000",
    600 => "00111110101000111011010001010000",
    601 => "00111110110010111110001101010000",
    602 => "00111110101000111011010001010000",
    603 => "00111110110010111110001101010000",
    604 => "00111110101000111011010001010000",
    605 => "00111110110010111110001101010000",
    606 => "00111111100000111101010110010110",
    607 => "00111110101000011110100010011011",
    608 => "00111110110011000001010011110111",
    609 => "00111110101000111011010100000110",
    610 => "00111110110010111110001101000010",
    611 => "00111110101000111011010001010000",
    612 => "00111110110010111110001101010001",
    613 => "00111110101000111011010001010000",
    614 => "00111110110010111110001101010001",
    615 => "00111110101000111011010001010000",
    616 => "00111110110010111110001101010001",
    617 => "00111111100000111101010110010110",
    618 => "00111110101000011110100010011011",
    619 => "00111111000001001111101110110100",
    620 => "00111110101001001010011110010010",
    621 => "00111111000001000000100101100000",
    622 => "00111110101001001010000001011110",
    623 => "00111111000001000000101101100101",
    624 => "00111110101001001010000001101101",
    625 => "00111111000001000000101101100011",
    626 => "00111110101001001010000001101101",
    627 => "00111111000001000000101101100011",
    628 => "00111111100010100110101101110000",
    629 => "00111110101000011110100010011011",
    630 => "00111110101011110011111110110000",
    631 => "00111110101000110101111000100011",
    632 => "00111110101011110011111001111011",
    633 => "00111110101000110101111000100001",
    634 => "00111110101011110011111001111011",
    635 => "00111110101000110101111000100001",
    636 => "00111110101011110011111001111011",
    637 => "00111110101000110101111000100001",
    638 => "00111110101011110011111001111011",
    639 => "00111111100000010011010100110101",
    640 => "00111110101000011110100010011011",
    641 => "00111111010100111001000101000010",
    642 => "00111110101001100101100001111011",
    643 => "00111111010010110010110001000000",
    644 => "00111110101001100011100001111100",
    645 => "00111111010010110101101011011100",
    646 => "00111110101001100011100100110101",
    647 => "00111111010010110101100111001011",
    648 => "00111110101001100011100100110001",
    649 => "00111111010010110101100111011001",
    650 => "00111111100111101010100000100110",
    651 => "00111110101000011110100010011011",
    652 => "00111110101000110100111001000100",
    653 => "00111110101000110100111010110000",
    654 => "00111110101000110100111010110000",
    655 => "00111110101000110100111010110000",
    656 => "00111110101000110100111010110000",
    657 => "00111110101000110100111010110000",
    658 => "00111110101000110100111010110000",
    659 => "00111110101000110100111010110000",
    660 => "00111110101000110100111010110000",
    661 => "00111111100000000011100011010000",
    662 => "00111110101000011110100010011011",
    663 => "00111110101000110100111001000100",
    664 => "00111110101011110011111001110011",
    665 => "00111110101000110101111000100001",
    666 => "00111110101011110011111001111011",
    667 => "00111110101000110101111000100001",
    668 => "00111110101011110011111001111011",
    669 => "00111110101000110101111000100001",
    670 => "00111110101011110011111001111011",
    671 => "00111110101000110101111000100001",
    672 => "00111111100000010011010100110101",
    673 => "00111110101000011110100010011011",
    674 => "00111111010100111000110000011011",
    675 => "00111110110001111100011100101001",
    676 => "00111111010001100100101101101001",
    677 => "00111110110001100101000001011000",
    678 => "00111111010001011011010011110110",
    679 => "00111110110001100011111001011000",
    680 => "00111111010001011010110111101011",
    681 => "00111110110001100011110110000001",
    682 => "00111111010001011010110110011001",
    683 => "00111111100111110010100101111011",
    684 => "00111110101000011110100010011011",
    685 => "00111110101011110011111110101111",
    686 => "00111110101011111010110111010000",
    687 => "00111110101011111011010100001101",
    688 => "00111110101011111011010110001001",
    689 => "00111110101011111011010110010001",
    690 => "00111110101011111011010110010010",
    691 => "00111110101011111011010110010010",
    692 => "00111110101011111011010110010010",
    693 => "00111110101011111011010110010010",
    694 => "00111111100000100100000101010100",
    695 => "00111110101000011110100010011011",
    696 => "00111111000001001111101110100011",
    697 => "00111110101110101011011011001101",
    698 => "00111111000001001000011000101000",
    699 => "00111110101110101001100111101110",
    700 => "00111111000001001000000000110000",
    701 => "00111110101110101001100001110111",
    702 => "00111111000001000111111111100010",
    703 => "00111110101110101001100001100011",
    704 => "00111111000001000111111111011110",
    705 => "00111111100011000100001000010100",
    706 => "00111110101000011110100010011011",
    707 => "00111110110011000001010011110110",
    708 => "00111110101100101001111100110011",
    709 => "00111110110011001110010110010101",
    710 => "00111110101100101011100101101101",
    711 => "00111110110011001110101001010110",
    712 => "00111110101100101011101000000111",
    713 => "00111110110011001110101001110000",
    714 => "00111110101100101011101000001010",
    715 => "00111110110011001110101001110001",
    716 => "00111111100001010010010110010001",
    717 => "00111110101000011110100010011011",
    718 => "00111110110011000001010011110111",
    719 => "00111110101100101001111100110100",
    720 => "00111110110011001110010110010110",
    721 => "00111110101100101011100101101101",
    722 => "00111110110011001110101001010111",
    723 => "00111110101100101011101000000111",
    724 => "00111110110011001110101001110010",
    725 => "00111110101100101011101000001001",
    726 => "00111110110011001110101001110011",
    727 => "00111111100001010010010110010010",
    728 => "00111110101000011110100010011011",
    729 => "00111111000001001111101110110100",
    730 => "00111110101110101011011011010010",
    731 => "00111111000001001000011000101000",
    732 => "00111110101110101001100111101110",
    733 => "00111111000001001000000000101110",
    734 => "00111110101110101001100001110110",
    735 => "00111111000001000111111111100001",
    736 => "00111110101110101001100001100010",
    737 => "00111111000001000111111111011100",
    738 => "00111111100011000100001000010011",
    739 => "00111110101000011110100010011011",
    740 => "00111110101011110011111110110000",
    741 => "00111110101011111010110111010000",
    742 => "00111110101011111011010100001110",
    743 => "00111110101011111011010110001001",
    744 => "00111110101011111011010110010010",
    745 => "00111110101011111011010110010010",
    746 => "00111110101011111011010110010010",
    747 => "00111110101011111011010110010010",
    748 => "00111110101011111011010110010010",
    749 => "00111111100000100100000101010100",
    750 => "00111110101000011110100010011011",
    751 => "00111111010100111001000101000010",
    752 => "00111110110001111100011110110001",
    753 => "00111111010001100100110011110111",
    754 => "00111110110001100101000010000111",
    755 => "00111111010001011011011001100011",
    756 => "00111110110001100011111010000101",
    757 => "00111111010001011010111101011000",
    758 => "00111110110001100011110110101100",
    759 => "00111111010001011010111100000101",
    760 => "00111111100111110010100111101111",
    761 => "00111110101000011110100010011011",
    762 => "00111110101000110100111001000100",
    763 => "00111110101011110011111001110011",
    764 => "00111110101000110101111000100001",
    765 => "00111110101011110011111001111011",
    766 => "00111110101000110101111000100001",
    767 => "00111110101011110011111001111011",
    768 => "00111110101000110101111000100001",
    769 => "00111110101011110011111001111011",
    770 => "00111110101000110101111000100001",
    771 => "00111111100000010011010100110101",
    772 => "00111110101000011110100010011011",
    773 => "00111110101000110100111001000100",
    774 => "00111110110010111110110001010100",
    775 => "00111110101000111011010001110001",
    776 => "00111110110010111110001101001101",
    777 => "00111110101000111011010001010000",
    778 => "00111110110010111110001101010000",
    779 => "00111110101000111011010001010000",
    780 => "00111110110010111110001101010000",
    781 => "00111110101000111011010001010000",
    782 => "00111111100000111101010110010110",
    783 => "00111110101000011110100010011011",
    784 => "00111111010100111000110000011111",
    785 => "00111111000000100101001011010001",
    786 => "00111111011000001010110100111110",
    787 => "00111111000000110111011011111110",
    788 => "00111111011000010110000110111100",
    789 => "00111111000000111000010100111101",
    790 => "00111111011000010110101001100000",
    791 => "00111111000000111000010111101010",
    792 => "00111111011000010110101011001010",
    793 => "00111111101011011001100000101001",
    794 => "00111110101000011110100010011011",
    795 => "00111110101011110011111110101111",
    796 => "00111110110011000101101100000111",
    797 => "00111110101100101010011111111110",
    798 => "00111110110011001110011100101100",
    799 => "00111110101100101011100110100000",
    800 => "00111110110011001110101001100000",
    801 => "00111110101100101011101000001000",
    802 => "00111110110011001110101001110000",
    803 => "00111110101100101011101000001010",
    804 => "00111111100001010010010110010001",
    805 => "00111110101000011110100010011011",
    806 => "00111111000001001111101110100011",
    807 => "00111110111010001001010000001001",
    808 => "00111111000100100011101110111010",
    809 => "00111110111011111101000001001010",
    810 => "00111111000101000111000101010100",
    811 => "00111110111100001110010110101110",
    812 => "00111111000101001100010000001011",
    813 => "00111110111100010000110110000110",
    814 => "00111111000101001100111111100001",
    815 => "00111111100101010100000000101111",
    816 => "00111110101000011110100010011011",
    817 => "00111110110011000001010011110110",
    818 => "00111110110100111110001110100110",
    819 => "00111110110101101000101010110011",
    820 => "00111110110101110111011001001001",
    821 => "00111110110101111100100001100010",
    822 => "00111110110101111110010100000101",
    823 => "00111110110101111110111100000100",
    824 => "00111110110101111111001010000001",
    825 => "00111110110101111111001110110111",
    826 => "00111111100010011001110001001010",
    827 => "00111110101000011110100010011011",
    828 => "00111110110011000001010011110111",
    829 => "00111110110100111110001110100111",
    830 => "00111110110101101000101010110100",
    831 => "00111110110101110111011001001001",
    832 => "00111110110101111100100001100011",
    833 => "00111110110101111110010100000110",
    834 => "00111110110101111110111100000101",
    835 => "00111110110101111111001010000000",
    836 => "00111110110101111111001110111001",
    837 => "00111111100010011001110001001011",
    838 => "00111110101000011110100010011011",
    839 => "00111111000001001111101110110100",
    840 => "00111110111010001001010000010100",
    841 => "00111111000100100011101110111100",
    842 => "00111110111011111101000001001100",
    843 => "00111111000101000111000101001111",
    844 => "00111110111100001110010110101110",
    845 => "00111111000101001100010000000110",
    846 => "00111110111100010000110110000011",
    847 => "00111111000101001100111111011010",
    848 => "00111111100101010100000000101101",
    849 => "00111110101000011110100010011011",
    850 => "00111110101011110011111110110000",
    851 => "00111110110011000101101100000111",
    852 => "00111110101100101010011111111110",
    853 => "00111110110011001110011100101100",
    854 => "00111110101100101011100110100000",
    855 => "00111110110011001110101001100000",
    856 => "00111110101100101011101000001000",
    857 => "00111110110011001110101001110000",
    858 => "00111110101100101011101000001010",
    859 => "00111111100001010010010110010010",
    860 => "00111110101000011110100010011011",
    861 => "00111111010100111001000101000010",
    862 => "00111111000000100101001101010000",
    863 => "00111111011000001010111001011010",
    864 => "00111111000000110111011100010100",
    865 => "00111111011000010110001010010110",
    866 => "00111111000000111000010101001110",
    867 => "00111111011000010110101100110001",
    868 => "00111111000000111000010111111010",
    869 => "00111111011000010110101110011001",
    870 => "00111111101011011001100001110000",
    871 => "00111110101000011110100010011011",
    872 => "00111110101000110100111001000100",
    873 => "00111110110010111110110001010100",
    874 => "00111110101000111011010001110001",
    875 => "00111110110010111110001101001101",
    876 => "00111110101000111011010001010000",
    877 => "00111110110010111110001101010000",
    878 => "00111110101000111011010001010000",
    879 => "00111110110010111110001101010000",
    880 => "00111110101000111011010001010000",
    881 => "00111111100000111101010110010110",
    882 => "00111110101000011110100010011011",
    883 => "00111110101000110100111001000100",
    884 => "00111111000001000111010010100010",
    885 => "00111110101001001010001110010000",
    886 => "00111111000001000000101001111111",
    887 => "00111110101001001010000001100111",
    888 => "00111111000001000000101101100011",
    889 => "00111110101001001010000001101110",
    890 => "00111111000001000000101101100010",
    891 => "00111110101001001010000001101110",
    892 => "00111111100010100110101101110000",
    893 => "00111110101000011110100010011011",
    894 => "00111111010100111000110000011011",
    895 => "00111111001011100001101100011011",
    896 => "00111111011011001111011100001111",
    897 => "00111111001011111101110101000010",
    898 => "00111111011011010000110000000110",
    899 => "00111111001011111101111001100011",
    900 => "00111111011011010000110000010010",
    901 => "00111111001011111101111001100010",
    902 => "00111111011011010000110000011000",
    903 => "00111111101110101100100000101110",
    904 => "00111110101000011110100010011011",
    905 => "00111110101011110011111110101111",
    906 => "00111111000000101111101111111011",
    907 => "00111110101110100011100001000101",
    908 => "00111111000001000110110000111101",
    909 => "00111110101110101001001110001100",
    910 => "00111111000001000111111011011101",
    911 => "00111110101110101001100000100010",
    912 => "00111111000001000111111111010000",
    913 => "00111110101110101001100001011110",
    914 => "00111111100011000100001000010011",
    915 => "00111110101000011110100010011011",
    916 => "00111111000001001111101110100011",
    917 => "00111111000110111000111010111111",
    918 => "00111111001001000110000000011010",
    919 => "00111111001001101100111100001111",
    920 => "00111111001001110110011001101011",
    921 => "00111111001001111000100111110100",
    922 => "00111111001001111001001000111101",
    923 => "00111111001001111001010000100100",
    924 => "00111111001001111001010010011010",
    925 => "00111111101001001100010011100000",
    926 => "00111110101000011110100010011011",
    927 => "00111110110011000001010011110110",
    928 => "00111111000010010010100110111000",
    929 => "00111110111010101111111110100110",
    930 => "00111111000100101111101101011110",
    931 => "00111110111100000010111101000010",
    932 => "00111111000101001000110110110000",
    933 => "00111110111100001111001101011110",
    934 => "00111111000101001100100000010111",
    935 => "00111110111100010000111101111001",
    936 => "00111111100101010011111111110010",
    937 => "00111110101000011110100010011011",
    938 => "00111110110011000001010011110111",
    939 => "00111111000010010010100110111001",
    940 => "00111110111010101111111110101001",
    941 => "00111111000100101111101101011110",
    942 => "00111110111100000010111101000110",
    943 => "00111111000101001000110110110010",
    944 => "00111110111100001111001101100010",
    945 => "00111111000101001100100000011001",
    946 => "00111110111100010000111101111101",
    947 => "00111111100101010011111111110011",
    948 => "00111110101000011110100010011011",
    949 => "00111111000001001111101110110100",
    950 => "00111111000110111000111011001001",
    951 => "00111111001001000110000000011110",
    952 => "00111111001001101100111100001101",
    953 => "00111111001001110110011001101001",
    954 => "00111111001001111000100111110010",
    955 => "00111111001001111001001000111010",
    956 => "00111111001001111001010000100101",
    957 => "00111111001001111001010010010111",
    958 => "00111111101001001100010011100000",
    959 => "00111110101000011110100010011011",
    960 => "00111110101011110011111110110000",
    961 => "00111111000000101111101111111100",
    962 => "00111110101110100011100001000110",
    963 => "00111111000001000110110000111101",
    964 => "00111110101110101001001110001100",
    965 => "00111111000001000111111011011101",
    966 => "00111110101110101001100000100010",
    967 => "00111111000001000111111111010000",
    968 => "00111110101110101001100001011111",
    969 => "00111111100011000100001000010011",
    970 => "00111110101000011110100010011011",
    971 => "00111111010100111001000101000010",
    972 => "00111111001011100001101110010001",
    973 => "00111111011011001111011100111100",
    974 => "00111111001011111101110101000111",
    975 => "00111111011011010000110000101100",
    976 => "00111111001011111101111001100100",
    977 => "00111111011011010000110000110110",
    978 => "00111111001011111101111001100100",
    979 => "00111111011011010000110000110110",
    980 => "00111111101110101100100000111000",
    981 => "00111110101000011110100010011011",
    982 => "00111110101000110100111001000100",
    983 => "00111111000001000111010010100010",
    984 => "00111110101001001010001110010000",
    985 => "00111111000001000000101001111111",
    986 => "00111110101001001010000001100111",
    987 => "00111111000001000000101101100011",
    988 => "00111110101001001010000001101110",
    989 => "00111111000001000000101101100010",
    990 => "00111110101001001010000001101110",
    991 => "00111111100010100110101101110000",
    992 => "00111110101000011110100010011011",
    993 => "00111110101000110100111001000100",
    994 => "00111111010100000111001100011000",
    995 => "00111110101001100100110011101010",
    996 => "00111111010010110011110011111111",
    997 => "00111110101001100011100010111110",
    998 => "00111111010010110101101010000000",
    999 => "00111110101001100011100100110011");

  component fsqrt is
    port (A : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          Q : out std_logic_vector (31 downto 0));
  end component fsqrt;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (3 downto 0) of std_logic_vector (31 downto 0);
  signal cc : buff := (others => (others => '0'));
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0'); 
  signal Q_buff : std_logic_vector (7 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
  signal i_isRunning : std_logic := 'U';
  signal i_result : std_logic := '1';
begin  -- architecture fsqrt_tb

  i_fsqrt : fsqrt port map (s_a,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk,Q_buff) is
    variable ss : character;
    variable count : integer := 4;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      case state is
        when "00" =>
          state <= "01";
        when "01" =>
          state <= "10";
        when "10" =>
          state <= "11";
        when others =>
          state <= "00";
      end case;
      s_a <= a_lut (addr);
      cc (conv_integer (state)) <= ans_lut (addr);
--      ccc <= cc ;

      if i_isRunning = '1' then  -- rising clock edge
        if cc (conv_integer (state)) = c and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 5 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;

  end process ram_loop;

end architecture;
