library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity finv is
  port (
    A : in std_logic_vector (31 downto 0);
    CLK : in std_logic;
    Q : out std_logic_vector (31 downto 0));
end entity finv;

architecture rtl of finv is

  function table(index: std_logic_vector(11 downto 0))
    return std_logic_vector
  is
    variable r : std_logic_vector(34 downto 0);
  begin
    case conv_integer(index) is
      when    0 => r := "11111111111010000000000000000000000";
      when    1 => r := "11111111111001111111111100000000001";
      when    2 => r := "11111111101001111111111000000000010";
      when    3 => r := "11111111101001111111110100000000101";
      when    4 => r := "11111111011001111111110000000001000";
      when    5 => r := "11111111011001111111101100000001101";
      when    6 => r := "11111111001001111111101000000010010";
      when    7 => r := "11111111001001111111100100000011001";
      when    8 => r := "11111110111001111111100000000100000";
      when    9 => r := "11111110111001111111011100000101001";
      when   10 => r := "11111110101001111111011000000110010";
      when   11 => r := "11111110101001111111010100000111101";
      when   12 => r := "11111110011001111111010000001001000";
      when   13 => r := "11111110011001111111001100001010101";
      when   14 => r := "11111110001001111111001000001100000";
      when   15 => r := "11111110001001111111000100001101111";
      when   16 => r := "11111101111001111111000000001111111";
      when   17 => r := "11111101111001111110111100010010000";
      when   18 => r := "11111101101001111110111000010100001";
      when   19 => r := "11111101101001111110110100010110100";
      when   20 => r := "11111101011001111110110000011000110";
      when   21 => r := "11111101011001111110101100011011011";
      when   22 => r := "11111101001001111110101000011110001";
      when   23 => r := "11111101001001111110100100100001000";
      when   24 => r := "11111100111001111110100000100011111";
      when   25 => r := "11111100111001111110011100100111000";
      when   26 => r := "11111100101001111110011000101001111";
      when   27 => r := "11111100101001111110010100101101010";
      when   28 => r := "11111100011001111110010000110000101";
      when   29 => r := "11111100011001111110001100110100010";
      when   30 => r := "11111100001001111110001000110111110";
      when   31 => r := "11111100001001111110000100111011101";
      when   32 => r := "11111011111001111110000000111111100";
      when   33 => r := "11111011111001111101111101000011101";
      when   34 => r := "11111011101001111101111001000111011";
      when   35 => r := "11111011101001111101110101001011110";
      when   36 => r := "11111011011001111101110001010000011";
      when   37 => r := "11111011011001111101101101010100111";
      when   38 => r := "11111011001101111101101001011001011";
      when   39 => r := "11111011001101111101100101011110001";
      when   40 => r := "11111010111101111101100001100011001";
      when   41 => r := "11111010111101111101011101101000010";
      when   42 => r := "11111010101101111101011001101101001";
      when   43 => r := "11111010101101111101010101110010100";
      when   44 => r := "11111010011101111101010001110111110";
      when   45 => r := "11111010011101111101001101111101010";
      when   46 => r := "11111010001101111101001010000010110";
      when   47 => r := "11111010001101111101000110001000101";
      when   48 => r := "11111001111101111101000010001110011";
      when   49 => r := "11111001111101111100111110010100011";
      when   50 => r := "11111001101101111100111010011010011";
      when   51 => r := "11111001101101111100110110100000101";
      when   52 => r := "11111001100001111100110010100111000";
      when   53 => r := "11111001100001111100101110101101100";
      when   54 => r := "11111001010001111100101010110011110";
      when   55 => r := "11111001010001111100100110111010100";
      when   56 => r := "11111001000001111100100011000001100";
      when   57 => r := "11111001000001111100011111001000011";
      when   58 => r := "11111000110001111100011011001111010";
      when   59 => r := "11111000110001111100010111010110100";
      when   60 => r := "11111000100001111100010011011101111";
      when   61 => r := "11111000100001111100001111100101011";
      when   62 => r := "11111000010001111100001011101100110";
      when   63 => r := "11111000010001111100000111110100100";
      when   64 => r := "11111000000101111100000011111100001";
      when   65 => r := "11111000000101111100000000000100000";
      when   66 => r := "11110111110101111011111100001011111";
      when   67 => r := "11110111110101111011111000010100000";
      when   68 => r := "11110111100101111011110100011100010";
      when   69 => r := "11110111100101111011110000100100101";
      when   70 => r := "11110111010101111011101100101101001";
      when   71 => r := "11110111010101111011101000110101110";
      when   72 => r := "11110111000101111011100100111110100";
      when   73 => r := "11110111000101111011100001000111011";
      when   74 => r := "11110110111001111011011101010000001";
      when   75 => r := "11110110111001111011011001011001010";
      when   76 => r := "11110110101001111011010101100010010";
      when   77 => r := "11110110101001111011010001101011101";
      when   78 => r := "11110110011001111011001101110101001";
      when   79 => r := "11110110011001111011001001111110110";
      when   80 => r := "11110110001001111011000110001000011";
      when   81 => r := "11110110001001111011000010010010010";
      when   82 => r := "11110101111001111010111110011100000";
      when   83 => r := "11110101111001111010111010100110001";
      when   84 => r := "11110101101101111010110110110000001";
      when   85 => r := "11110101101101111010110010111010100";
      when   86 => r := "11110101011101111010101111000100101";
      when   87 => r := "11110101011101111010101011001111001";
      when   88 => r := "11110101001101111010100111011001110";
      when   89 => r := "11110101001101111010100011100100100";
      when   90 => r := "11110100111101111010011111101111010";
      when   91 => r := "11110100111101111010011011111010010";
      when   92 => r := "11110100110001111010011000000101100";
      when   93 => r := "11110100110001111010010100010000110";
      when   94 => r := "11110100100001111010010000011100000";
      when   95 => r := "11110100100001111010001100100111011";
      when   96 => r := "11110100010001111010001000110010111";
      when   97 => r := "11110100010001111010000100111110101";
      when   98 => r := "11110100000001111010000001001010001";
      when   99 => r := "11110100000001111001111101010110001";
      when  100 => r := "11110011110101111001111001100010001";
      when  101 => r := "11110011110101111001110101101110011";
      when  102 => r := "11110011100101111001110001111010011";
      when  103 => r := "11110011100101111001101110000110111";
      when  104 => r := "11110011010101111001101010010011000";
      when  105 => r := "11110011010101111001100110011111110";
      when  106 => r := "11110011001001111001100010101100100";
      when  107 => r := "11110011001001111001011110111001011";
      when  108 => r := "11110010111001111001011011000110001";
      when  109 => r := "11110010111001111001010111010011010";
      when  110 => r := "11110010101001111001010011100000100";
      when  111 => r := "11110010101001111001001111101101111";
      when  112 => r := "11110010011101111001001011111011000";
      when  113 => r := "11110010011101111001001000001000100";
      when  114 => r := "11110010001101111001000100010110001";
      when  115 => r := "11110010001101111001000000100100000";
      when  116 => r := "11110001111101111000111100110001111";
      when  117 => r := "11110001111101111000111000111111111";
      when  118 => r := "11110001101101111000110101001101110";
      when  119 => r := "11110001101101111000110001011100000";
      when  120 => r := "11110001100001111000101101101010011";
      when  121 => r := "11110001100001111000101001111000111";
      when  122 => r := "11110001010001111000100110000111010";
      when  123 => r := "11110001010001111000100010010110000";
      when  124 => r := "11110001000001111000011110100100111";
      when  125 => r := "11110001000001111000011010110011111";
      when  126 => r := "11110000110101111000010111000010101";
      when  127 => r := "11110000110101111000010011010001111";
      when  128 => r := "11110000100101111000001111100000111";
      when  129 => r := "11110000100101111000001011110000010";
      when  130 => r := "11110000011001111000000111111111110";
      when  131 => r := "11110000011001111000000100001111011";
      when  132 => r := "11110000001001111000000000011110111";
      when  133 => r := "11110000001001110111111100101110110";
      when  134 => r := "11101111111001110111111000111110101";
      when  135 => r := "11101111111001110111110101001110110";
      when  136 => r := "11101111101101110111110001011110110";
      when  137 => r := "11101111101101110111101101101111001";
      when  138 => r := "11101111011101110111101001111111100";
      when  139 => r := "11101111011101110111100110010000000";
      when  140 => r := "11101111001101110111100010100000100";
      when  141 => r := "11101111001101110111011110110001010";
      when  142 => r := "11101111000001110111011011000001111";
      when  143 => r := "11101111000001110111010111010010111";
      when  144 => r := "11101110110001110111010011100100000";
      when  145 => r := "11101110110001110111001111110101010";
      when  146 => r := "11101110100101110111001100000110100";
      when  147 => r := "11101110100101110111001000010111111";
      when  148 => r := "11101110010101110111000100101001010";
      when  149 => r := "11101110010101110111000000111010111";
      when  150 => r := "11101110000101110110111101001100100";
      when  151 => r := "11101110000101110110111001011110100";
      when  152 => r := "11101101111001110110110101110000010";
      when  153 => r := "11101101111001110110110010000010011";
      when  154 => r := "11101101101001110110101110010100100";
      when  155 => r := "11101101101001110110101010100110111";
      when  156 => r := "11101101011101110110100110111001001";
      when  157 => r := "11101101011101110110100011001011110";
      when  158 => r := "11101101001101110110011111011110010";
      when  159 => r := "11101101001101110110011011110001001";
      when  160 => r := "11101101000001110110011000000011111";
      when  161 => r := "11101101000001110110010100010110111";
      when  162 => r := "11101100110001110110010000101001110";
      when  163 => r := "11101100110001110110001100111101000";
      when  164 => r := "11101100100001110110001001010000010";
      when  165 => r := "11101100100001110110000101100011110";
      when  166 => r := "11101100010101110110000001110111010";
      when  167 => r := "11101100010101110101111110001010111";
      when  168 => r := "11101100000101110101111010011110011";
      when  169 => r := "11101100000101110101110110110010010";
      when  170 => r := "11101011111001110101110011000110010";
      when  171 => r := "11101011111001110101101111011010011";
      when  172 => r := "11101011101001110101101011101110100";
      when  173 => r := "11101011101001110101101000000010111";
      when  174 => r := "11101011011101110101100100010111010";
      when  175 => r := "11101011011101110101100000101011110";
      when  176 => r := "11101011001101110101011101000000010";
      when  177 => r := "11101011001101110101011001010101000";
      when  178 => r := "11101011000001110101010101101001110";
      when  179 => r := "11101011000001110101010001111110110";
      when  180 => r := "11101010110001110101001110010011110";
      when  181 => r := "11101010110001110101001010101000111";
      when  182 => r := "11101010100101110101000110111110010";
      when  183 => r := "11101010100101110101000011010011101";
      when  184 => r := "11101010010101110100111111101001000";
      when  185 => r := "11101010010101110100111011111110110";
      when  186 => r := "11101010001001110100111000010100011";
      when  187 => r := "11101010001001110100110100101010010";
      when  188 => r := "11101001111001110100110001000000001";
      when  189 => r := "11101001111001110100101101010110010";
      when  190 => r := "11101001101101110100101001101100001";
      when  191 => r := "11101001101101110100100110000010100";
      when  192 => r := "11101001011101110100100010011000111";
      when  193 => r := "11101001011101110100011110101111011";
      when  194 => r := "11101001010001110100011011000101111";
      when  195 => r := "11101001010001110100010111011100101";
      when  196 => r := "11101001000001110100010011110011011";
      when  197 => r := "11101001000001110100010000001010011";
      when  198 => r := "11101000110101110100001100100001010";
      when  199 => r := "11101000110101110100001000111000011";
      when  200 => r := "11101000100101110100000101001111110";
      when  201 => r := "11101000100101110100000001100111001";
      when  202 => r := "11101000011001110011111101111110011";
      when  203 => r := "11101000011001110011111010010110000";
      when  204 => r := "11101000001001110011110110101101101";
      when  205 => r := "11101000001001110011110011000101100";
      when  206 => r := "11100111111101110011101111011101010";
      when  207 => r := "11100111111101110011101011110101011";
      when  208 => r := "11100111101101110011101000001101010";
      when  209 => r := "11100111101101110011100100100101101";
      when  210 => r := "11100111100001110011100000111101111";
      when  211 => r := "11100111100001110011011101010110011";
      when  212 => r := "11100111010101110011011001101110101";
      when  213 => r := "11100111010101110011010110000111010";
      when  214 => r := "11100111000101110011010010100000010";
      when  215 => r := "11100111000101110011001110111001001";
      when  216 => r := "11100110111001110011001011010010000";
      when  217 => r := "11100110111001110011000111101011001";
      when  218 => r := "11100110101001110011000100000100000";
      when  219 => r := "11100110101001110011000000011101011";
      when  220 => r := "11100110011101110010111100110110110";
      when  221 => r := "11100110011101110010111001010000010";
      when  222 => r := "11100110001101110010110101101001111";
      when  223 => r := "11100110001101110010110010000011101";
      when  224 => r := "11100110000001110010101110011101010";
      when  225 => r := "11100110000001110010101010110111010";
      when  226 => r := "11100101110101110010100111010001011";
      when  227 => r := "11100101110101110010100011101011101";
      when  228 => r := "11100101100101110010100000000101101";
      when  229 => r := "11100101100101110010011100100000001";
      when  230 => r := "11100101011001110010011000111010011";
      when  231 => r := "11100101011001110010010101010100111";
      when  232 => r := "11100101001001110010010001101111101";
      when  233 => r := "11100101001001110010001110001010011";
      when  234 => r := "11100100111101110010001010100101010";
      when  235 => r := "11100100111101110010000111000000011";
      when  236 => r := "11100100110001110010000011011011010";
      when  237 => r := "11100100110001110001111111110110100";
      when  238 => r := "11100100100001110001111100010001111";
      when  239 => r := "11100100100001110001111000101101011";
      when  240 => r := "11100100010101110001110101001000110";
      when  241 => r := "11100100010101110001110001100100011";
      when  242 => r := "11100100001001110001101110000000001";
      when  243 => r := "11100100001001110001101010011100000";
      when  244 => r := "11100011111001110001100110110111101";
      when  245 => r := "11100011111001110001100011010011110";
      when  246 => r := "11100011101101110001011111110000001";
      when  247 => r := "11100011101101110001011100001100011";
      when  248 => r := "11100011011101110001011000101000100";
      when  249 => r := "11100011011101110001010101000101000";
      when  250 => r := "11100011010001110001010001100001101";
      when  251 => r := "11100011010001110001001101111110011";
      when  252 => r := "11100011000101110001001010011010110";
      when  253 => r := "11100011000101110001000110110111110";
      when  254 => r := "11100010110101110001000011010100111";
      when  255 => r := "11100010110101110000111111110010000";
      when  256 => r := "11100010101001110000111100001111000";
      when  257 => r := "11100010101001110000111000101100011";
      when  258 => r := "11100010011101110000110101001001111";
      when  259 => r := "11100010011101110000110001100111011";
      when  260 => r := "11100010001101110000101110000100111";
      when  261 => r := "11100010001101110000101010100010101";
      when  262 => r := "11100010000001110000100111000000011";
      when  263 => r := "11100010000001110000100011011110011";
      when  264 => r := "11100001110101110000011111111100010";
      when  265 => r := "11100001110101110000011100011010100";
      when  266 => r := "11100001101001110000011000111000101";
      when  267 => r := "11100001101001110000010101010111000";
      when  268 => r := "11100001011001110000010001110101010";
      when  269 => r := "11100001011001110000001110010011111";
      when  270 => r := "11100001001101110000001010110010011";
      when  271 => r := "11100001001101110000000111010001010";
      when  272 => r := "11100001000001110000000011110000001";
      when  273 => r := "11100001000001110000000000001111000";
      when  274 => r := "11100000110001101111111100101110001";
      when  275 => r := "11100000110001101111111001001101011";
      when  276 => r := "11100000100101101111110101101100100";
      when  277 => r := "11100000100101101111110010001011111";
      when  278 => r := "11100000011001101111101110101011010";
      when  279 => r := "11100000011001101111101011001010111";
      when  280 => r := "11100000001001101111100111101010100";
      when  281 => r := "11100000001001101111100100001010011";
      when  282 => r := "11011111111101101111100000101010001";
      when  283 => r := "11011111111101101111011101001010001";
      when  284 => r := "11011111110001101111011001101010001";
      when  285 => r := "11011111110001101111010110001010011";
      when  286 => r := "11011111100101101111010010101010100";
      when  287 => r := "11011111100101101111001111001011000";
      when  288 => r := "11011111010101101111001011101011011";
      when  289 => r := "11011111010101101111001000001100001";
      when  290 => r := "11011111001001101111000100101100101";
      when  291 => r := "11011111001001101111000001001101100";
      when  292 => r := "11011110111101101110111101101110010";
      when  293 => r := "11011110111101101110111010001111011";
      when  294 => r := "11011110110001101110110110110000100";
      when  295 => r := "11011110110001101110110011010001101";
      when  296 => r := "11011110100001101110101111110010111";
      when  297 => r := "11011110100001101110101100010100011";
      when  298 => r := "11011110010101101110101000110101111";
      when  299 => r := "11011110010101101110100101010111100";
      when  300 => r := "11011110001001101110100001111001001";
      when  301 => r := "11011110001001101110011110011011000";
      when  302 => r := "11011101111101101110011010111100111";
      when  303 => r := "11011101111101101110010111011110111";
      when  304 => r := "11011101101101101110010100000000111";
      when  305 => r := "11011101101101101110010000100011001";
      when  306 => r := "11011101100001101110001101000101011";
      when  307 => r := "11011101100001101110001001100111111";
      when  308 => r := "11011101010101101110000110001010010";
      when  309 => r := "11011101010101101110000010101101000";
      when  310 => r := "11011101001001101101111111001111100";
      when  311 => r := "11011101001001101101111011110010011";
      when  312 => r := "11011100111101101101111000010101100";
      when  313 => r := "11011100111101101101110100111000100";
      when  314 => r := "11011100101101101101110001011011011";
      when  315 => r := "11011100101101101101101101111110101";
      when  316 => r := "11011100100001101101101010100010000";
      when  317 => r := "11011100100001101101100111000101100";
      when  318 => r := "11011100010101101101100011101000111";
      when  319 => r := "11011100010101101101100000001100100";
      when  320 => r := "11011100001001101101011100110000011";
      when  321 => r := "11011100001001101101011001010100010";
      when  322 => r := "11011011111101101101010101110111111";
      when  323 => r := "11011011111101101101010010011011111";
      when  324 => r := "11011011101101101101001111000000000";
      when  325 => r := "11011011101101101101001011100100010";
      when  326 => r := "11011011100001101101001000001000100";
      when  327 => r := "11011011100001101101000100101101000";
      when  328 => r := "11011011010101101101000001010001100";
      when  329 => r := "11011011010101101100111101110110001";
      when  330 => r := "11011011001001101100111010011010101";
      when  331 => r := "11011011001001101100110110111111100";
      when  332 => r := "11011010111101101100110011100100100";
      when  333 => r := "11011010111101101100110000001001100";
      when  334 => r := "11011010110001101100101100101110101";
      when  335 => r := "11011010110001101100101001010011111";
      when  336 => r := "11011010100001101100100101111000111";
      when  337 => r := "11011010100001101100100010011110011";
      when  338 => r := "11011010010101101100011111000100000";
      when  339 => r := "11011010010101101100011011101001110";
      when  340 => r := "11011010001001101100011000001111011";
      when  341 => r := "11011010001001101100010100110101010";
      when  342 => r := "11011001111101101100010001011010111";
      when  343 => r := "11011001111101101100001110000001000";
      when  344 => r := "11011001110001101100001010100110111";
      when  345 => r := "11011001110001101100000111001101000";
      when  346 => r := "11011001100101101100000011110011100";
      when  347 => r := "11011001100101101100000000011001111";
      when  348 => r := "11011001011001101011111101000000010";
      when  349 => r := "11011001011001101011111001100110111";
      when  350 => r := "11011001001001101011110110001101100";
      when  351 => r := "11011001001001101011110010110100011";
      when  352 => r := "11011000111101101011101111011011010";
      when  353 => r := "11011000111101101011101100000010010";
      when  354 => r := "11011000110001101011101000101001010";
      when  355 => r := "11011000110001101011100101010000100";
      when  356 => r := "11011000100101101011100001110111101";
      when  357 => r := "11011000100101101011011110011111000";
      when  358 => r := "11011000011001101011011011000110100";
      when  359 => r := "11011000011001101011010111101110001";
      when  360 => r := "11011000001101101011010100010101100";
      when  361 => r := "11011000001101101011010000111101011";
      when  362 => r := "11011000000001101011001101100101001";
      when  363 => r := "11011000000001101011001010001101000";
      when  364 => r := "11010111110101101011000110110101010";
      when  365 => r := "11010111110101101011000011011101011";
      when  366 => r := "11010111101001101011000000000101100";
      when  367 => r := "11010111101001101010111100101101111";
      when  368 => r := "11010111011001101010111001010110010";
      when  369 => r := "11010111011001101010110101111110111";
      when  370 => r := "11010111001101101010110010100111010";
      when  371 => r := "11010111001101101010101111010000000";
      when  372 => r := "11010111000001101010101011111000111";
      when  373 => r := "11010111000001101010101000100001110";
      when  374 => r := "11010110110101101010100101001010110";
      when  375 => r := "11010110110101101010100001110100000";
      when  376 => r := "11010110101001101010011110011101001";
      when  377 => r := "11010110101001101010011011000110100";
      when  378 => r := "11010110011101101010010111101111110";
      when  379 => r := "11010110011101101010010100011001011";
      when  380 => r := "11010110010001101010010001000010110";
      when  381 => r := "11010110010001101010001101101100100";
      when  382 => r := "11010110000101101010001010010110001";
      when  383 => r := "11010110000101101010000111000000001";
      when  384 => r := "11010101111001101010000011101010000";
      when  385 => r := "11010101111001101010000000010100001";
      when  386 => r := "11010101101101101001111100111110010";
      when  387 => r := "11010101101101101001111001101000101";
      when  388 => r := "11010101100001101001110110010010111";
      when  389 => r := "11010101100001101001110010111101011";
      when  390 => r := "11010101010101101001101111100111111";
      when  391 => r := "11010101010101101001101100010010100";
      when  392 => r := "11010101001001101001101000111101010";
      when  393 => r := "11010101001001101001100101101000001";
      when  394 => r := "11010100111101101001100010010010111";
      when  395 => r := "11010100111101101001011110111101111";
      when  396 => r := "11010100110001101001011011101000111";
      when  397 => r := "11010100110001101001011000010100001";
      when  398 => r := "11010100100101101001010100111111011";
      when  399 => r := "11010100100101101001010001101010111";
      when  400 => r := "11010100011001101001001110010110010";
      when  401 => r := "11010100011001101001001011000001111";
      when  402 => r := "11010100001101101001000111101101100";
      when  403 => r := "11010100001101101001000100011001010";
      when  404 => r := "11010100000001101001000001000101001";
      when  405 => r := "11010100000001101000111101110001001";
      when  406 => r := "11010011110101101000111010011101010";
      when  407 => r := "11010011110101101000110111001001011";
      when  408 => r := "11010011101001101000110011110101100";
      when  409 => r := "11010011101001101000110000100001111";
      when  410 => r := "11010011011101101000101101001110010";
      when  411 => r := "11010011011101101000101001111010110";
      when  412 => r := "11010011010001101000100110100111100";
      when  413 => r := "11010011010001101000100011010100010";
      when  414 => r := "11010011000101101000100000000001000";
      when  415 => r := "11010011000101101000011100101101111";
      when  416 => r := "11010010111001101000011001011010110";
      when  417 => r := "11010010111001101000010110000111111";
      when  418 => r := "11010010101101101000010010110101001";
      when  419 => r := "11010010101101101000001111100010011";
      when  420 => r := "11010010100001101000001100001111100";
      when  421 => r := "11010010100001101000001000111101000";
      when  422 => r := "11010010010101101000000101101010110";
      when  423 => r := "11010010010101101000000010011000011";
      when  424 => r := "11010010001001100111111111000101111";
      when  425 => r := "11010010001001100111111011110011110";
      when  426 => r := "11010001111101100111111000100001101";
      when  427 => r := "11010001111101100111110101001111101";
      when  428 => r := "11010001110001100111110001111101111";
      when  429 => r := "11010001110001100111101110101100001";
      when  430 => r := "11010001100101100111101011011010010";
      when  431 => r := "11010001100101100111101000001000110";
      when  432 => r := "11010001011001100111100100110111001";
      when  433 => r := "11010001011001100111100001100101110";
      when  434 => r := "11010001001101100111011110010100010";
      when  435 => r := "11010001001101100111011011000011001";
      when  436 => r := "11010001000001100111010111110001111";
      when  437 => r := "11010001000001100111010100100000111";
      when  438 => r := "11010000110101100111010001010000000";
      when  439 => r := "11010000110101100111001101111111001";
      when  440 => r := "11010000101001100111001010101110001";
      when  441 => r := "11010000101001100111000111011101100";
      when  442 => r := "11010000011101100111000100001100111";
      when  443 => r := "11010000011101100111000000111100100";
      when  444 => r := "11010000010001100110111101101100000";
      when  445 => r := "11010000010001100110111010011011110";
      when  446 => r := "11010000000101100110110111001011100";
      when  447 => r := "11010000000101100110110011111011011";
      when  448 => r := "11001111111001100110110000101011010";
      when  449 => r := "11001111111001100110101101011011011";
      when  450 => r := "11001111101101100110101010001011101";
      when  451 => r := "11001111101101100110100110111011111";
      when  452 => r := "11001111100001100110100011101100000";
      when  453 => r := "11001111100001100110100000011100100";
      when  454 => r := "11001111010101100110011101001100110";
      when  455 => r := "11001111010101100110011001111101011";
      when  456 => r := "11001111001101100110010110101110001";
      when  457 => r := "11001111001101100110010011011111000";
      when  458 => r := "11001111000001100110010000001111101";
      when  459 => r := "11001111000001100110001101000000101";
      when  460 => r := "11001110110101100110001001110001101";
      when  461 => r := "11001110110101100110000110100010110";
      when  462 => r := "11001110101001100110000011010011111";
      when  463 => r := "11001110101001100110000000000101010";
      when  464 => r := "11001110011101100101111100110110110";
      when  465 => r := "11001110011101100101111001101000011";
      when  466 => r := "11001110010001100101110110011001101";
      when  467 => r := "11001110010001100101110011001011011";
      when  468 => r := "11001110000101100101101111111101010";
      when  469 => r := "11001110000101100101101100101111001";
      when  470 => r := "11001101111001100101101001100001001";
      when  471 => r := "11001101111001100101100110010011010";
      when  472 => r := "11001101101101100101100011000101010";
      when  473 => r := "11001101101101100101011111110111100";
      when  474 => r := "11001101100001100101011100101001110";
      when  475 => r := "11001101100001100101011001011100001";
      when  476 => r := "11001101011001100101010110001110101";
      when  477 => r := "11001101011001100101010011000001010";
      when  478 => r := "11001101001101100101001111110011111";
      when  479 => r := "11001101001101100101001100100110110";
      when  480 => r := "11001101000001100101001001011001011";
      when  481 => r := "11001101000001100101000110001100011";
      when  482 => r := "11001100110101100101000010111111011";
      when  483 => r := "11001100110101100100111111110010101";
      when  484 => r := "11001100101001100100111100100101110";
      when  485 => r := "11001100101001100100111001011001001";
      when  486 => r := "11001100011101100100110110001100100";
      when  487 => r := "11001100011101100100110011000000001";
      when  488 => r := "11001100010001100100101111110011011";
      when  489 => r := "11001100010001100100101100100111000";
      when  490 => r := "11001100001001100100101001011010111";
      when  491 => r := "11001100001001100100100110001110110";
      when  492 => r := "11001011111101100100100011000010101";
      when  493 => r := "11001011111101100100011111110110110";
      when  494 => r := "11001011110001100100011100101010110";
      when  495 => r := "11001011110001100100011001011110111";
      when  496 => r := "11001011100101100100010110010011001";
      when  497 => r := "11001011100101100100010011000111101";
      when  498 => r := "11001011011001100100001111111100000";
      when  499 => r := "11001011011001100100001100110000101";
      when  500 => r := "11001011001101100100001001100101010";
      when  501 => r := "11001011001101100100000110011010000";
      when  502 => r := "11001011000101100100000011001110110";
      when  503 => r := "11001011000101100100000000000011101";
      when  504 => r := "11001010111001100011111100111000100";
      when  505 => r := "11001010111001100011111001101101101";
      when  506 => r := "11001010101101100011110110100010110";
      when  507 => r := "11001010101101100011110011011000001";
      when  508 => r := "11001010100001100011110000001101011";
      when  509 => r := "11001010100001100011101101000010111";
      when  510 => r := "11001010010101100011101001111000011";
      when  511 => r := "11001010010101100011100110101110000";
      when  512 => r := "11001010001001100011100011100011011";
      when  513 => r := "11001010001001100011100000011001010";
      when  514 => r := "11001010000001100011011101001111010";
      when  515 => r := "11001010000001100011011010000101001";
      when  516 => r := "11001001110101100011010110111011010";
      when  517 => r := "11001001110101100011010011110001011";
      when  518 => r := "11001001101001100011010000100111100";
      when  519 => r := "11001001101001100011001101011101111";
      when  520 => r := "11001001011101100011001010010100001";
      when  521 => r := "11001001011101100011000111001010110";
      when  522 => r := "11001001010001100011000100000001001";
      when  523 => r := "11001001010001100011000000110111111";
      when  524 => r := "11001001001001100010111101101110101";
      when  525 => r := "11001001001001100010111010100101011";
      when  526 => r := "11001000111101100010110111011100010";
      when  527 => r := "11001000111101100010110100010011011";
      when  528 => r := "11001000110001100010110001001010011";
      when  529 => r := "11001000110001100010101110000001101";
      when  530 => r := "11001000100101100010101010111000110";
      when  531 => r := "11001000100101100010100111110000010";
      when  532 => r := "11001000011101100010100100100111101";
      when  533 => r := "11001000011101100010100001011111010";
      when  534 => r := "11001000010001100010011110010110111";
      when  535 => r := "11001000010001100010011011001110100";
      when  536 => r := "11001000000101100010011000000110010";
      when  537 => r := "11001000000101100010010100111110010";
      when  538 => r := "11000111111001100010010001110110000";
      when  539 => r := "11000111111001100010001110101110000";
      when  540 => r := "11000111101101100010001011100110001";
      when  541 => r := "11000111101101100010001000011110011";
      when  542 => r := "11000111100101100010000101010110101";
      when  543 => r := "11000111100101100010000010001111000";
      when  544 => r := "11000111011001100001111111000111101";
      when  545 => r := "11000111011001100001111100000000001";
      when  546 => r := "11000111001101100001111000111000110";
      when  547 => r := "11000111001101100001110101110001101";
      when  548 => r := "11000111000001100001110010101010010";
      when  549 => r := "11000111000001100001101111100011010";
      when  550 => r := "11000110111001100001101100011100000";
      when  551 => r := "11000110111001100001101001010101001";
      when  552 => r := "11000110101101100001100110001110011";
      when  553 => r := "11000110101101100001100011000111110";
      when  554 => r := "11000110100001100001100000000000110";
      when  555 => r := "11000110100001100001011100111010010";
      when  556 => r := "11000110011001100001011001110011110";
      when  557 => r := "11000110011001100001010110101101011";
      when  558 => r := "11000110001101100001010011100111001";
      when  559 => r := "11000110001101100001010000100001000";
      when  560 => r := "11000110000001100001001101011010101";
      when  561 => r := "11000110000001100001001010010100100";
      when  562 => r := "11000101110101100001000111001110100";
      when  563 => r := "11000101110101100001000100001000101";
      when  564 => r := "11000101101101100001000001000010111";
      when  565 => r := "11000101101101100000111101111101001";
      when  566 => r := "11000101100001100000111010110111011";
      when  567 => r := "11000101100001100000110111110001111";
      when  568 => r := "11000101010101100000110100101100011";
      when  569 => r := "11000101010101100000110001100111000";
      when  570 => r := "11000101001101100000101110100001101";
      when  571 => r := "11000101001101100000101011011100011";
      when  572 => r := "11000101000001100000101000010111001";
      when  573 => r := "11000101000001100000100101010010001";
      when  574 => r := "11000100110101100000100010001101010";
      when  575 => r := "11000100110101100000011111001000011";
      when  576 => r := "11000100101001100000011100000011100";
      when  577 => r := "11000100101001100000011000111110111";
      when  578 => r := "11000100100001100000010101111010001";
      when  579 => r := "11000100100001100000010010110101101";
      when  580 => r := "11000100010101100000001111110001001";
      when  581 => r := "11000100010101100000001100101100110";
      when  582 => r := "11000100001001100000001001101000011";
      when  583 => r := "11000100001001100000000110100100010";
      when  584 => r := "11000100000001100000000011100000000";
      when  585 => r := "11000100000001100000000000011011111";
      when  586 => r := "11000011110101011111111101011000000";
      when  587 => r := "11000011110101011111111010010100010";
      when  588 => r := "11000011101001011111110111010000010";
      when  589 => r := "11000011101001011111110100001100101";
      when  590 => r := "11000011100001011111110001001001000";
      when  591 => r := "11000011100001011111101110000101100";
      when  592 => r := "11000011010101011111101011000010000";
      when  593 => r := "11000011010101011111100111111110101";
      when  594 => r := "11000011001001011111100100111011011";
      when  595 => r := "11000011001001011111100001111000001";
      when  596 => r := "11000011000001011111011110110101000";
      when  597 => r := "11000011000001011111011011110010000";
      when  598 => r := "11000010110101011111011000101110111";
      when  599 => r := "11000010110101011111010101101100001";
      when  600 => r := "11000010101001011111010010101001001";
      when  601 => r := "11000010101001011111001111100110100";
      when  602 => r := "11000010100001011111001100100011111";
      when  603 => r := "11000010100001011111001001100001011";
      when  604 => r := "11000010010101011111000110011110111";
      when  605 => r := "11000010010101011111000011011100100";
      when  606 => r := "11000010001001011111000000011010000";
      when  607 => r := "11000010001001011110111101010111111";
      when  608 => r := "11000010000001011110111010010101110";
      when  609 => r := "11000010000001011110110111010011110";
      when  610 => r := "11000001110101011110110100010001110";
      when  611 => r := "11000001110101011110110001001111111";
      when  612 => r := "11000001101101011110101110001110000";
      when  613 => r := "11000001101101011110101011001100011";
      when  614 => r := "11000001100001011110101000001010110";
      when  615 => r := "11000001100001011110100101001001010";
      when  616 => r := "11000001010101011110100010000111101";
      when  617 => r := "11000001010101011110011111000110010";
      when  618 => r := "11000001001101011110011100000100110";
      when  619 => r := "11000001001101011110011001000011101";
      when  620 => r := "11000001000001011110010110000010011";
      when  621 => r := "11000001000001011110010011000001011";
      when  622 => r := "11000000110101011110010000000000100";
      when  623 => r := "11000000110101011110001100111111110";
      when  624 => r := "11000000101101011110001001111110101";
      when  625 => r := "11000000101101011110000110111101111";
      when  626 => r := "11000000100001011110000011111101001";
      when  627 => r := "11000000100001011110000000111100101";
      when  628 => r := "11000000011001011101111101111100010";
      when  629 => r := "11000000011001011101111010111011111";
      when  630 => r := "11000000001101011101110111111011011";
      when  631 => r := "11000000001101011101110100111011001";
      when  632 => r := "11000000000001011101110001111011001";
      when  633 => r := "11000000000001011101101110111011001";
      when  634 => r := "10111111111001011101101011111010111";
      when  635 => r := "10111111111001011101101000111011000";
      when  636 => r := "10111111101101011101100101111011000";
      when  637 => r := "10111111101101011101100010111011011";
      when  638 => r := "10111111100101011101011111111011110";
      when  639 => r := "10111111100101011101011100111100001";
      when  640 => r := "10111111011001011101011001111100100";
      when  641 => r := "10111111011001011101010110111101001";
      when  642 => r := "10111111001101011101010011111101110";
      when  643 => r := "10111111001101011101010000111110100";
      when  644 => r := "10111111000101011101001101111111011";
      when  645 => r := "10111111000101011101001011000000010";
      when  646 => r := "10111110111001011101001000000001000";
      when  647 => r := "10111110111001011101000101000010001";
      when  648 => r := "10111110110001011101000010000011001";
      when  649 => r := "10111110110001011100111111000100011";
      when  650 => r := "10111110100101011100111100000101101";
      when  651 => r := "10111110100101011100111001000111000";
      when  652 => r := "10111110011101011100110110001000100";
      when  653 => r := "10111110011101011100110011001010000";
      when  654 => r := "10111110010001011100110000001011100";
      when  655 => r := "10111110010001011100101101001101010";
      when  656 => r := "10111110000101011100101010001111001";
      when  657 => r := "10111110000101011100100111010001001";
      when  658 => r := "10111101111101011100100100010010111";
      when  659 => r := "10111101111101011100100001010100111";
      when  660 => r := "10111101110001011100011110010111000";
      when  661 => r := "10111101110001011100011011011001001";
      when  662 => r := "10111101101001011100011000011011011";
      when  663 => r := "10111101101001011100010101011101110";
      when  664 => r := "10111101011101011100010010100000000";
      when  665 => r := "10111101011101011100001111100010101";
      when  666 => r := "10111101010101011100001100100100111";
      when  667 => r := "10111101010101011100001001100111101";
      when  668 => r := "10111101001001011100000110101010011";
      when  669 => r := "10111101001001011100000011101101010";
      when  670 => r := "10111101000001011100000000110000010";
      when  671 => r := "10111101000001011011111101110011010";
      when  672 => r := "10111100110101011011111010110110000";
      when  673 => r := "10111100110101011011110111111001010";
      when  674 => r := "10111100101001011011110100111100011";
      when  675 => r := "10111100101001011011110001111111110";
      when  676 => r := "10111100100001011011101111000011001";
      when  677 => r := "10111100100001011011101100000110101";
      when  678 => r := "10111100010101011011101001001010001";
      when  679 => r := "10111100010101011011100110001101110";
      when  680 => r := "10111100001101011011100011010001001";
      when  681 => r := "10111100001101011011100000010101000";
      when  682 => r := "10111100000001011011011101011000110";
      when  683 => r := "10111100000001011011011010011100110";
      when  684 => r := "10111011111001011011010111100000110";
      when  685 => r := "10111011111001011011010100100100110";
      when  686 => r := "10111011101101011011010001101000110";
      when  687 => r := "10111011101101011011001110101101001";
      when  688 => r := "10111011100101011011001011110001011";
      when  689 => r := "10111011100101011011001000110101110";
      when  690 => r := "10111011011001011011000101111010001";
      when  691 => r := "10111011011001011011000010111110110";
      when  692 => r := "10111011010001011011000000000011011";
      when  693 => r := "10111011010001011010111101001000001";
      when  694 => r := "10111011000101011010111010001100110";
      when  695 => r := "10111011000101011010110111010001101";
      when  696 => r := "10111010111101011010110100010110110";
      when  697 => r := "10111010111101011010110001011011110";
      when  698 => r := "10111010110001011010101110100000110";
      when  699 => r := "10111010110001011010101011100110000";
      when  700 => r := "10111010101001011010101000101011001";
      when  701 => r := "10111010101001011010100101110000100";
      when  702 => r := "10111010011101011010100010110101110";
      when  703 => r := "10111010011101011010011111111011011";
      when  704 => r := "10111010010101011010011101000000101";
      when  705 => r := "10111010010101011010011010000110011";
      when  706 => r := "10111010001001011010010111001100010";
      when  707 => r := "10111010001001011010010100010010001";
      when  708 => r := "10111010000001011010010001010111111";
      when  709 => r := "10111010000001011010001110011101111";
      when  710 => r := "10111001110101011010001011100011110";
      when  711 => r := "10111001110101011010001000101001111";
      when  712 => r := "10111001101101011010000101101111111";
      when  713 => r := "10111001101101011010000010110110001";
      when  714 => r := "10111001100001011001111111111100101";
      when  715 => r := "10111001100001011001111101000011001";
      when  716 => r := "10111001011001011001111010001001100";
      when  717 => r := "10111001011001011001110111010000001";
      when  718 => r := "10111001010001011001110100010110101";
      when  719 => r := "10111001010001011001110001011101011";
      when  720 => r := "10111001000101011001101110100100010";
      when  721 => r := "10111001000101011001101011101011001";
      when  722 => r := "10111000111101011001101000110010000";
      when  723 => r := "10111000111101011001100101111001000";
      when  724 => r := "10111000110001011001100011000000000";
      when  725 => r := "10111000110001011001100000000111010";
      when  726 => r := "10111000101001011001011101001110100";
      when  727 => r := "10111000101001011001011010010101111";
      when  728 => r := "10111000011101011001010111011101010";
      when  729 => r := "10111000011101011001010100100100110";
      when  730 => r := "10111000010101011001010001101100010";
      when  731 => r := "10111000010101011001001110110011111";
      when  732 => r := "10111000001001011001001011111011011";
      when  733 => r := "10111000001001011001001001000011010";
      when  734 => r := "10111000000001011001000110001011010";
      when  735 => r := "10111000000001011001000011010011010";
      when  736 => r := "10110111111001011001000000011011001";
      when  737 => r := "10110111111001011000111101100011010";
      when  738 => r := "10110111101101011000111010101011010";
      when  739 => r := "10110111101101011000110111110011101";
      when  740 => r := "10110111100101011000110100111011111";
      when  741 => r := "10110111100101011000110010000100010";
      when  742 => r := "10110111011001011000101111001100101";
      when  743 => r := "10110111011001011000101100010101010";
      when  744 => r := "10110111010001011000101001011110000";
      when  745 => r := "10110111010001011000100110100110101";
      when  746 => r := "10110111000101011000100011101111011";
      when  747 => r := "10110111000101011000100000111000011";
      when  748 => r := "10110110111101011000011110000001001";
      when  749 => r := "10110110111101011000011011001010001";
      when  750 => r := "10110110110101011000011000010011001";
      when  751 => r := "10110110110101011000010101011100011";
      when  752 => r := "10110110101001011000010010100101101";
      when  753 => r := "10110110101001011000001111101111000";
      when  754 => r := "10110110100001011000001100111000010";
      when  755 => r := "10110110100001011000001010000001110";
      when  756 => r := "10110110010101011000000111001011010";
      when  757 => r := "10110110010101011000000100010100111";
      when  758 => r := "10110110001101011000000001011110100";
      when  759 => r := "10110110001101010111111110101000010";
      when  760 => r := "10110110000101010111111011110010000";
      when  761 => r := "10110110000101010111111000111100000";
      when  762 => r := "10110101111001010111110110000110000";
      when  763 => r := "10110101111001010111110011010000001";
      when  764 => r := "10110101110001010111110000011010001";
      when  765 => r := "10110101110001010111101101100100011";
      when  766 => r := "10110101100101010111101010101110100";
      when  767 => r := "10110101100101010111100111111001000";
      when  768 => r := "10110101011101010111100101000011011";
      when  769 => r := "10110101011101010111100010001101111";
      when  770 => r := "10110101010101010111011111011000100";
      when  771 => r := "10110101010101010111011100100011001";
      when  772 => r := "10110101001001010111011001101101101";
      when  773 => r := "10110101001001010111010110111000100";
      when  774 => r := "10110101000001010111010100000011100";
      when  775 => r := "10110101000001010111010001001110100";
      when  776 => r := "10110100110101010111001110011001101";
      when  777 => r := "10110100110101010111001011100100110";
      when  778 => r := "10110100101101010111001000101111101";
      when  779 => r := "10110100101101010111000101111010111";
      when  780 => r := "10110100100101010111000011000110001";
      when  781 => r := "10110100100101010111000000010001101";
      when  782 => r := "10110100011001010110111101011101001";
      when  783 => r := "10110100011001010110111010101000110";
      when  784 => r := "10110100010001010110110111110100010";
      when  785 => r := "10110100010001010110110100111111111";
      when  786 => r := "10110100001001010110110010001011101";
      when  787 => r := "10110100001001010110101111010111100";
      when  788 => r := "10110011111101010110101100100011100";
      when  789 => r := "10110011111101010110101001101111100";
      when  790 => r := "10110011110101010110100110111011101";
      when  791 => r := "10110011110101010110100100000111110";
      when  792 => r := "10110011101101010110100001010011110";
      when  793 => r := "10110011101101010110011110100000001";
      when  794 => r := "10110011100001010110011011101100100";
      when  795 => r := "10110011100001010110011000111001000";
      when  796 => r := "10110011011001010110010110000101001";
      when  797 => r := "10110011011001010110010011010001110";
      when  798 => r := "10110011001101010110010000011110100";
      when  799 => r := "10110011001101010110001101101011010";
      when  800 => r := "10110011000101010110001010111000000";
      when  801 => r := "10110011000101010110001000000101000";
      when  802 => r := "10110010111101010110000101010010000";
      when  803 => r := "10110010111101010110000010011111000";
      when  804 => r := "10110010110001010101111111101100000";
      when  805 => r := "10110010110001010101111100111001001";
      when  806 => r := "10110010101001010101111010000110011";
      when  807 => r := "10110010101001010101110111010011110";
      when  808 => r := "10110010100001010101110100100001000";
      when  809 => r := "10110010100001010101110001101110011";
      when  810 => r := "10110010010101010101101110111011111";
      when  811 => r := "10110010010101010101101100001001100";
      when  812 => r := "10110010001101010101101001010111010";
      when  813 => r := "10110010001101010101100110100101001";
      when  814 => r := "10110010000101010101100011110010110";
      when  815 => r := "10110010000101010101100001000000101";
      when  816 => r := "10110001111001010101011110001110101";
      when  817 => r := "10110001111001010101011011011100110";
      when  818 => r := "10110001110001010101011000101010110";
      when  819 => r := "10110001110001010101010101111001000";
      when  820 => r := "10110001101001010101010011000111000";
      when  821 => r := "10110001101001010101010000010101011";
      when  822 => r := "10110001100001010101001101100011110";
      when  823 => r := "10110001100001010101001010110010010";
      when  824 => r := "10110001010101010101001000000000111";
      when  825 => r := "10110001010101010101000101001111101";
      when  826 => r := "10110001001101010101000010011110001";
      when  827 => r := "10110001001101010100111111101100111";
      when  828 => r := "10110001000101010100111100111011110";
      when  829 => r := "10110001000101010100111010001010101";
      when  830 => r := "10110000111001010100110111011001100";
      when  831 => r := "10110000111001010100110100101000101";
      when  832 => r := "10110000110001010100110001110111101";
      when  833 => r := "10110000110001010100101111000110111";
      when  834 => r := "10110000101001010100101100010110000";
      when  835 => r := "10110000101001010100101001100101011";
      when  836 => r := "10110000011101010100100110110100110";
      when  837 => r := "10110000011101010100100100000100010";
      when  838 => r := "10110000010101010100100001010011110";
      when  839 => r := "10110000010101010100011110100011100";
      when  840 => r := "10110000001101010100011011110011001";
      when  841 => r := "10110000001101010100011001000011000";
      when  842 => r := "10110000000101010100010110010010110";
      when  843 => r := "10110000000101010100010011100010110";
      when  844 => r := "10101111111001010100010000110010100";
      when  845 => r := "10101111111001010100001110000010101";
      when  846 => r := "10101111110001010100001011010010101";
      when  847 => r := "10101111110001010100001000100010111";
      when  848 => r := "10101111101001010100000101110011010";
      when  849 => r := "10101111101001010100000011000011101";
      when  850 => r := "10101111011101010100000000010011111";
      when  851 => r := "10101111011101010011111101100100011";
      when  852 => r := "10101111010101010011111010110101000";
      when  853 => r := "10101111010101010011111000000101101";
      when  854 => r := "10101111001101010011110101010110010";
      when  855 => r := "10101111001101010011110010100111000";
      when  856 => r := "10101111000101010011101111110111101";
      when  857 => r := "10101111000101010011101101001000101";
      when  858 => r := "10101110111001010011101010011001100";
      when  859 => r := "10101110111001010011100111101010101";
      when  860 => r := "10101110110001010011100100111011101";
      when  861 => r := "10101110110001010011100010001100111";
      when  862 => r := "10101110101001010011011111011110010";
      when  863 => r := "10101110101001010011011100101111100";
      when  864 => r := "10101110100001010011011010000000111";
      when  865 => r := "10101110100001010011010111010010011";
      when  866 => r := "10101110010101010011010100100011110";
      when  867 => r := "10101110010101010011010001110101100";
      when  868 => r := "10101110001101010011001111000111000";
      when  869 => r := "10101110001101010011001100011000111";
      when  870 => r := "10101110000101010011001001101010101";
      when  871 => r := "10101110000101010011000110111100101";
      when  872 => r := "10101101111101010011000100001110011";
      when  873 => r := "10101101111101010011000001100000011";
      when  874 => r := "10101101110001010010111110110010101";
      when  875 => r := "10101101110001010010111100000100110";
      when  876 => r := "10101101101001010010111001010110111";
      when  877 => r := "10101101101001010010110110101001010";
      when  878 => r := "10101101100001010010110011111011100";
      when  879 => r := "10101101100001010010110001001101111";
      when  880 => r := "10101101011001010010101110100000011";
      when  881 => r := "10101101011001010010101011110011000";
      when  882 => r := "10101101010001010010101001000101110";
      when  883 => r := "10101101010001010010100110011000100";
      when  884 => r := "10101101000101010010100011101011010";
      when  885 => r := "10101101000101010010100000111110001";
      when  886 => r := "10101100111101010010011110010000111";
      when  887 => r := "10101100111101010010011011100100000";
      when  888 => r := "10101100110101010010011000110111001";
      when  889 => r := "10101100110101010010010110001010010";
      when  890 => r := "10101100101101010010010011011101011";
      when  891 => r := "10101100101101010010010000110000110";
      when  892 => r := "10101100100001010010001110000100000";
      when  893 => r := "10101100100001010010001011010111100";
      when  894 => r := "10101100011001010010001000101010111";
      when  895 => r := "10101100011001010010000101111110100";
      when  896 => r := "10101100010001010010000011010001111";
      when  897 => r := "10101100010001010010000000100101101";
      when  898 => r := "10101100001001010001111101111001101";
      when  899 => r := "10101100001001010001111011001101011";
      when  900 => r := "10101100000001010001111000100001010";
      when  901 => r := "10101100000001010001110101110101010";
      when  902 => r := "10101011110101010001110011001001001";
      when  903 => r := "10101011110101010001110000011101010";
      when  904 => r := "10101011101101010001101101110001011";
      when  905 => r := "10101011101101010001101011000101110";
      when  906 => r := "10101011100101010001101000011001111";
      when  907 => r := "10101011100101010001100101101110011";
      when  908 => r := "10101011011101010001100011000010111";
      when  909 => r := "10101011011101010001100000010111011";
      when  910 => r := "10101011010101010001011101101011111";
      when  911 => r := "10101011010101010001011011000000101";
      when  912 => r := "10101011001001010001011000010101011";
      when  913 => r := "10101011001001010001010101101010010";
      when  914 => r := "10101011000001010001010010111110111";
      when  915 => r := "10101011000001010001010000010011111";
      when  916 => r := "10101010111001010001001101101000111";
      when  917 => r := "10101010111001010001001010111110000";
      when  918 => r := "10101010110001010001001000010011000";
      when  919 => r := "10101010110001010001000101101000001";
      when  920 => r := "10101010101001010001000010111101100";
      when  921 => r := "10101010101001010001000000010010111";
      when  922 => r := "10101010100001010000111101101000001";
      when  923 => r := "10101010100001010000111010111101101";
      when  924 => r := "10101010010101010000111000010011001";
      when  925 => r := "10101010010101010000110101101000110";
      when  926 => r := "10101010001101010000110010111110011";
      when  927 => r := "10101010001101010000110000010100010";
      when  928 => r := "10101010000101010000101101101010000";
      when  929 => r := "10101010000101010000101010111111111";
      when  930 => r := "10101001111101010000101000010101111";
      when  931 => r := "10101001111101010000100101101011111";
      when  932 => r := "10101001110101010000100011000001111";
      when  933 => r := "10101001110101010000100000011000000";
      when  934 => r := "10101001101101010000011101101110010";
      when  935 => r := "10101001101101010000011011000100100";
      when  936 => r := "10101001100001010000011000011010111";
      when  937 => r := "10101001100001010000010101110001011";
      when  938 => r := "10101001011001010000010011000111111";
      when  939 => r := "10101001011001010000010000011110100";
      when  940 => r := "10101001010001010000001101110100111";
      when  941 => r := "10101001010001010000001011001011101";
      when  942 => r := "10101001001001010000001000100010010";
      when  943 => r := "10101001001001010000000101111001000";
      when  944 => r := "10101001000001010000000011010000001";
      when  945 => r := "10101001000001010000000000100111000";
      when  946 => r := "10101000111001001111111101111101111";
      when  947 => r := "10101000111001001111111011010101000";
      when  948 => r := "10101000101101001111111000101100010";
      when  949 => r := "10101000101101001111110110000011100";
      when  950 => r := "10101000100101001111110011011010101";
      when  951 => r := "10101000100101001111110000110010000";
      when  952 => r := "10101000011101001111101110001001101";
      when  953 => r := "10101000011101001111101011100001001";
      when  954 => r := "10101000010101001111101000111000101";
      when  955 => r := "10101000010101001111100110010000010";
      when  956 => r := "10101000001101001111100011100111110";
      when  957 => r := "10101000001101001111100000111111101";
      when  958 => r := "10101000000101001111011110010111100";
      when  959 => r := "10101000000101001111011011101111011";
      when  960 => r := "10100111111101001111011001000111010";
      when  961 => r := "10100111111101001111010110011111010";
      when  962 => r := "10100111110101001111010011110111010";
      when  963 => r := "10100111110101001111010001001111100";
      when  964 => r := "10100111101001001111001110100111110";
      when  965 => r := "10100111101001001111001100000000000";
      when  966 => r := "10100111100001001111001001011000100";
      when  967 => r := "10100111100001001111000110110001000";
      when  968 => r := "10100111011001001111000100001001011";
      when  969 => r := "10100111011001001111000001100001111";
      when  970 => r := "10100111010001001110111110111010011";
      when  971 => r := "10100111010001001110111100010011001";
      when  972 => r := "10100111001001001110111001101011110";
      when  973 => r := "10100111001001001110110111000100101";
      when  974 => r := "10100111000001001110110100011101101";
      when  975 => r := "10100111000001001110110001110110100";
      when  976 => r := "10100110111001001110101111001111100";
      when  977 => r := "10100110111001001110101100101000101";
      when  978 => r := "10100110110001001110101010000001111";
      when  979 => r := "10100110110001001110100111011011001";
      when  980 => r := "10100110101001001110100100110100011";
      when  981 => r := "10100110101001001110100010001101110";
      when  982 => r := "10100110011101001110011111100110111";
      when  983 => r := "10100110011101001110011101000000011";
      when  984 => r := "10100110010101001110011010011010001";
      when  985 => r := "10100110010101001110010111110011110";
      when  986 => r := "10100110001101001110010101001101011";
      when  987 => r := "10100110001101001110010010100111001";
      when  988 => r := "10100110000101001110010000000000110";
      when  989 => r := "10100110000101001110001101011010110";
      when  990 => r := "10100101111101001110001010110100110";
      when  991 => r := "10100101111101001110001000001110111";
      when  992 => r := "10100101110101001110000101101000101";
      when  993 => r := "10100101110101001110000011000010110";
      when  994 => r := "10100101101101001110000000011100111";
      when  995 => r := "10100101101101001101111101110111010";
      when  996 => r := "10100101100101001101111011010001100";
      when  997 => r := "10100101100101001101111000101011111";
      when  998 => r := "10100101011101001101110110000110011";
      when  999 => r := "10100101011101001101110011100001000";
      when 1000 => r := "10100101010101001101110000111011011";
      when 1001 => r := "10100101010101001101101110010110000";
      when 1002 => r := "10100101001101001101101011110000101";
      when 1003 => r := "10100101001101001101101001001011100";
      when 1004 => r := "10100101000101001101100110100110100";
      when 1005 => r := "10100101000101001101100100000001011";
      when 1006 => r := "10100100111001001101100001011100010";
      when 1007 => r := "10100100111001001101011110110111011";
      when 1008 => r := "10100100110001001101011100010010011";
      when 1009 => r := "10100100110001001101011001101101101";
      when 1010 => r := "10100100101001001101010111001000110";
      when 1011 => r := "10100100101001001101010100100100001";
      when 1012 => r := "10100100100001001101010001111111100";
      when 1013 => r := "10100100100001001101001111011011000";
      when 1014 => r := "10100100011001001101001100110110100";
      when 1015 => r := "10100100011001001101001010010010000";
      when 1016 => r := "10100100010001001101000111101101101";
      when 1017 => r := "10100100010001001101000101001001011";
      when 1018 => r := "10100100001001001101000010100101000";
      when 1019 => r := "10100100001001001101000000000000111";
      when 1020 => r := "10100100000001001100111101011100110";
      when 1021 => r := "10100100000001001100111010111000110";
      when 1022 => r := "10100011111001001100111000010100101";
      when 1023 => r := "10100011111001001100110101110000101";
      when 1024 => r := "10100011110001001100110011001100110";
      when 1025 => r := "10100011110001001100110000101001000";
      when 1026 => r := "10100011101001001100101110000101001";
      when 1027 => r := "10100011101001001100101011100001100";
      when 1028 => r := "10100011100001001100101000111110000";
      when 1029 => r := "10100011100001001100100110011010011";
      when 1030 => r := "10100011011001001100100011110110111";
      when 1031 => r := "10100011011001001100100001010011100";
      when 1032 => r := "10100011010001001100011110110000001";
      when 1033 => r := "10100011010001001100011100001100111";
      when 1034 => r := "10100011001001001100011001101001101";
      when 1035 => r := "10100011001001001100010111000110100";
      when 1036 => r := "10100011000001001100010100100011010";
      when 1037 => r := "10100011000001001100010010000000010";
      when 1038 => r := "10100010111001001100001111011101010";
      when 1039 => r := "10100010111001001100001100111010011";
      when 1040 => r := "10100010110001001100001010010111100";
      when 1041 => r := "10100010110001001100000111110100110";
      when 1042 => r := "10100010101001001100000101010001111";
      when 1043 => r := "10100010101001001100000010101111010";
      when 1044 => r := "10100010100001001100000000001100110";
      when 1045 => r := "10100010100001001011111101101010010";
      when 1046 => r := "10100010011001001011111011000111110";
      when 1047 => r := "10100010011001001011111000100101011";
      when 1048 => r := "10100010010001001011110110000010111";
      when 1049 => r := "10100010010001001011110011100000101";
      when 1050 => r := "10100010001001001011110000111110100";
      when 1051 => r := "10100010001001001011101110011100011";
      when 1052 => r := "10100001111101001011101011111010010";
      when 1053 => r := "10100001111101001011101001011000011";
      when 1054 => r := "10100001110101001011100110110110001";
      when 1055 => r := "10100001110101001011100100010100010";
      when 1056 => r := "10100001101101001011100001110010100";
      when 1057 => r := "10100001101101001011011111010000111";
      when 1058 => r := "10100001100101001011011100101111000";
      when 1059 => r := "10100001100101001011011010001101011";
      when 1060 => r := "10100001011101001011010111101011110";
      when 1061 => r := "10100001011101001011010101001010010";
      when 1062 => r := "10100001010101001011010010101000110";
      when 1063 => r := "10100001010101001011010000000111011";
      when 1064 => r := "10100001001101001011001101100110000";
      when 1065 => r := "10100001001101001011001011000100110";
      when 1066 => r := "10100001000101001011001000100011100";
      when 1067 => r := "10100001000101001011000110000010011";
      when 1068 => r := "10100000111101001011000011100001011";
      when 1069 => r := "10100000111101001011000001000000011";
      when 1070 => r := "10100000110101001010111110011111011";
      when 1071 => r := "10100000110101001010111011111110100";
      when 1072 => r := "10100000101101001010111001011101101";
      when 1073 => r := "10100000101101001010110110111100111";
      when 1074 => r := "10100000100101001010110100011100000";
      when 1075 => r := "10100000100101001010110001111011011";
      when 1076 => r := "10100000011101001010101111011010110";
      when 1077 => r := "10100000011101001010101100111010010";
      when 1078 => r := "10100000011001001010101010011001110";
      when 1079 => r := "10100000011001001010100111111001011";
      when 1080 => r := "10100000010001001010100101011001000";
      when 1081 => r := "10100000010001001010100010111000110";
      when 1082 => r := "10100000001001001010100000011000100";
      when 1083 => r := "10100000001001001010011101111000011";
      when 1084 => r := "10100000000001001010011011011000010";
      when 1085 => r := "10100000000001001010011000111000010";
      when 1086 => r := "10011111111001001010010110011000010";
      when 1087 => r := "10011111111001001010010011111000011";
      when 1088 => r := "10011111110001001010010001011000100";
      when 1089 => r := "10011111110001001010001110111000110";
      when 1090 => r := "10011111101001001010001100011001000";
      when 1091 => r := "10011111101001001010001001111001011";
      when 1092 => r := "10011111100001001010000111011001100";
      when 1093 => r := "10011111100001001010000100111010000";
      when 1094 => r := "10011111011001001010000010011010110";
      when 1095 => r := "10011111011001001001111111111011011";
      when 1096 => r := "10011111010001001001111101011100000";
      when 1097 => r := "10011111010001001001111010111100110";
      when 1098 => r := "10011111001001001001111000011101010";
      when 1099 => r := "10011111001001001001110101111110001";
      when 1100 => r := "10011111000001001001110011011111000";
      when 1101 => r := "10011111000001001001110001000000000";
      when 1102 => r := "10011110111001001001101110100001000";
      when 1103 => r := "10011110111001001001101100000010001";
      when 1104 => r := "10011110110001001001101001100011011";
      when 1105 => r := "10011110110001001001100111000100100";
      when 1106 => r := "10011110101001001001100100100101110";
      when 1107 => r := "10011110101001001001100010000111001";
      when 1108 => r := "10011110100001001001011111101000100";
      when 1109 => r := "10011110100001001001011101001010000";
      when 1110 => r := "10011110011001001001011010101011010";
      when 1111 => r := "10011110011001001001011000001100111";
      when 1112 => r := "10011110010001001001010101101110100";
      when 1113 => r := "10011110010001001001010011010000010";
      when 1114 => r := "10011110001001001001010000110001111";
      when 1115 => r := "10011110001001001001001110010011110";
      when 1116 => r := "10011110000001001001001011110101100";
      when 1117 => r := "10011110000001001001001001010111100";
      when 1118 => r := "10011101111001001001000110111001011";
      when 1119 => r := "10011101111001001001000100011011011";
      when 1120 => r := "10011101110001001001000001111101100";
      when 1121 => r := "10011101110001001000111111011111110";
      when 1122 => r := "10011101101001001000111101000010000";
      when 1123 => r := "10011101101001001000111010100100010";
      when 1124 => r := "10011101100001001000111000000110101";
      when 1125 => r := "10011101100001001000110101101001000";
      when 1126 => r := "10011101011101001000110011001011100";
      when 1127 => r := "10011101011101001000110000101110001";
      when 1128 => r := "10011101010101001000101110010000101";
      when 1129 => r := "10011101010101001000101011110011010";
      when 1130 => r := "10011101001101001000101001010110000";
      when 1131 => r := "10011101001101001000100110111000110";
      when 1132 => r := "10011101000101001000100100011011101";
      when 1133 => r := "10011101000101001000100001111110101";
      when 1134 => r := "10011100111101001000011111100001100";
      when 1135 => r := "10011100111101001000011101000100100";
      when 1136 => r := "10011100110101001000011010100111011";
      when 1137 => r := "10011100110101001000011000001010101";
      when 1138 => r := "10011100101101001000010101101101111";
      when 1139 => r := "10011100101101001000010011010001001";
      when 1140 => r := "10011100100101001000010000110100011";
      when 1141 => r := "10011100100101001000001110010111111";
      when 1142 => r := "10011100011101001000001011111011001";
      when 1143 => r := "10011100011101001000001001011110110";
      when 1144 => r := "10011100010101001000000111000010011";
      when 1145 => r := "10011100010101001000000100100110000";
      when 1146 => r := "10011100001101001000000010001001100";
      when 1147 => r := "10011100001101000111111111101101011";
      when 1148 => r := "10011100000101000111111101010001001";
      when 1149 => r := "10011100000101000111111010110101000";
      when 1150 => r := "10011100000001000111111000011000101";
      when 1151 => r := "10011100000001000111110101111100101";
      when 1152 => r := "10011011111001000111110011100000111";
      when 1153 => r := "10011011111001000111110001000101000";
      when 1154 => r := "10011011110001000111101110101001000";
      when 1155 => r := "10011011110001000111101100001101010";
      when 1156 => r := "10011011101001000111101001110001100";
      when 1157 => r := "10011011101001000111100111010101111";
      when 1158 => r := "10011011100001000111100100111010010";
      when 1159 => r := "10011011100001000111100010011110110";
      when 1160 => r := "10011011011001000111100000000011010";
      when 1161 => r := "10011011011001000111011101100111111";
      when 1162 => r := "10011011010001000111011011001100011";
      when 1163 => r := "10011011010001000111011000110001001";
      when 1164 => r := "10011011001001000111010110010101110";
      when 1165 => r := "10011011001001000111010011111010101";
      when 1166 => r := "10011011000001000111010001011111011";
      when 1167 => r := "10011011000001000111001111000100011";
      when 1168 => r := "10011010111101000111001100101001001";
      when 1169 => r := "10011010111101000111001010001110010";
      when 1170 => r := "10011010110101000111000111110011011";
      when 1171 => r := "10011010110101000111000101011000101";
      when 1172 => r := "10011010101101000111000010111101100";
      when 1173 => r := "10011010101101000111000000100010111";
      when 1174 => r := "10011010100101000110111110001000011";
      when 1175 => r := "10011010100101000110111011101101110";
      when 1176 => r := "10011010011101000110111001010011010";
      when 1177 => r := "10011010011101000110110110111000110";
      when 1178 => r := "10011010010101000110110100011110001";
      when 1179 => r := "10011010010101000110110010000011111";
      when 1180 => r := "10011010001101000110101111101001011";
      when 1181 => r := "10011010001101000110101101001111001";
      when 1182 => r := "10011010000101000110101010110101000";
      when 1183 => r := "10011010000101000110101000011010111";
      when 1184 => r := "10011010000001000110100110000000111";
      when 1185 => r := "10011010000001000110100011100110111";
      when 1186 => r := "10011001111001000110100001001100111";
      when 1187 => r := "10011001111001000110011110110011000";
      when 1188 => r := "10011001110001000110011100011000111";
      when 1189 => r := "10011001110001000110011001111111001";
      when 1190 => r := "10011001101001000110010111100101100";
      when 1191 => r := "10011001101001000110010101001011110";
      when 1192 => r := "10011001100001000110010010110010001";
      when 1193 => r := "10011001100001000110010000011000101";
      when 1194 => r := "10011001011001000110001101111111000";
      when 1195 => r := "10011001011001000110001011100101101";
      when 1196 => r := "10011001010001000110001001001100010";
      when 1197 => r := "10011001010001000110000110110011000";
      when 1198 => r := "10011001001101000110000100011001100";
      when 1199 => r := "10011001001101000110000010000000010";
      when 1200 => r := "10011001000101000101111111100111001";
      when 1201 => r := "10011001000101000101111101001110001";
      when 1202 => r := "10011000111101000101111010110101000";
      when 1203 => r := "10011000111101000101111000011100001";
      when 1204 => r := "10011000110101000101110110000011001";
      when 1205 => r := "10011000110101000101110011101010010";
      when 1206 => r := "10011000101101000101110001010001100";
      when 1207 => r := "10011000101101000101101110111000110";
      when 1208 => r := "10011000100101000101101100011111111";
      when 1209 => r := "10011000100101000101101010000111011";
      when 1210 => r := "10011000011101000101100111101110110";
      when 1211 => r := "10011000011101000101100101010110010";
      when 1212 => r := "10011000011001000101100010111110000";
      when 1213 => r := "10011000011001000101100000100101101";
      when 1214 => r := "10011000010001000101011110001101001";
      when 1215 => r := "10011000010001000101011011110100111";
      when 1216 => r := "10011000001001000101011001011100011";
      when 1217 => r := "10011000001001000101010111000100010";
      when 1218 => r := "10011000000001000101010100101100001";
      when 1219 => r := "10011000000001000101010010010100001";
      when 1220 => r := "10010111111001000101001111111100001";
      when 1221 => r := "10010111111001000101001101100100010";
      when 1222 => r := "10010111110001000101001011001100010";
      when 1223 => r := "10010111110001000101001000110100011";
      when 1224 => r := "10010111101101000101000110011100101";
      when 1225 => r := "10010111101101000101000100000100111";
      when 1226 => r := "10010111100101000101000001101101011";
      when 1227 => r := "10010111100101000100111111010101110";
      when 1228 => r := "10010111011101000100111100111110010";
      when 1229 => r := "10010111011101000100111010100110110";
      when 1230 => r := "10010111010101000100111000001111001";
      when 1231 => r := "10010111010101000100110101110111111";
      when 1232 => r := "10010111001101000100110011100000011";
      when 1233 => r := "10010111001101000100110001001001001";
      when 1234 => r := "10010111001001000100101110110010000";
      when 1235 => r := "10010111001001000100101100011010111";
      when 1236 => r := "10010111000001000100101010000011101";
      when 1237 => r := "10010111000001000100100111101100101";
      when 1238 => r := "10010110111001000100100101010101110";
      when 1239 => r := "10010110111001000100100010111110111";
      when 1240 => r := "10010110110001000100100000100111111";
      when 1241 => r := "10010110110001000100011110010001001";
      when 1242 => r := "10010110101001000100011011111010011";
      when 1243 => r := "10010110101001000100011001100011110";
      when 1244 => r := "10010110100001000100010111001100111";
      when 1245 => r := "10010110100001000100010100110110011";
      when 1246 => r := "10010110011101000100010010011111110";
      when 1247 => r := "10010110011101000100010000001001010";
      when 1248 => r := "10010110010101000100001101110011000";
      when 1249 => r := "10010110010101000100001011011100101";
      when 1250 => r := "10010110001101000100001001000110010";
      when 1251 => r := "10010110001101000100000110110000001";
      when 1252 => r := "10010110000101000100000100011001110";
      when 1253 => r := "10010110000101000100000010000011110";
      when 1254 => r := "10010101111101000011111111101101100";
      when 1255 => r := "10010101111101000011111101010111100";
      when 1256 => r := "10010101111001000011111011000001101";
      when 1257 => r := "10010101111001000011111000101011110";
      when 1258 => r := "10010101110001000011110110010101110";
      when 1259 => r := "10010101110001000011110100000000000";
      when 1260 => r := "10010101101001000011110001101010010";
      when 1261 => r := "10010101101001000011101111010100101";
      when 1262 => r := "10010101100001000011101100111110111";
      when 1263 => r := "10010101100001000011101010101001011";
      when 1264 => r := "10010101011101000011101000010011111";
      when 1265 => r := "10010101011101000011100101111110100";
      when 1266 => r := "10010101010101000011100011101000111";
      when 1267 => r := "10010101010101000011100001010011101";
      when 1268 => r := "10010101001101000011011110111110011";
      when 1269 => r := "10010101001101000011011100101001001";
      when 1270 => r := "10010101000101000011011010010011111";
      when 1271 => r := "10010101000101000011010111111110110";
      when 1272 => r := "10010100111101000011010101101001101";
      when 1273 => r := "10010100111101000011010011010100101";
      when 1274 => r := "10010100111001000011010000111111110";
      when 1275 => r := "10010100111001000011001110101010111";
      when 1276 => r := "10010100110001000011001100010110000";
      when 1277 => r := "10010100110001000011001010000001010";
      when 1278 => r := "10010100101001000011000111101100011";
      when 1279 => r := "10010100101001000011000101010111110";
      when 1280 => r := "10010100100001000011000011000011000";
      when 1281 => r := "10010100100001000011000000101110100";
      when 1282 => r := "10010100011101000010111110011010000";
      when 1283 => r := "10010100011101000010111100000101101";
      when 1284 => r := "10010100010101000010111001110001001";
      when 1285 => r := "10010100010101000010110111011100110";
      when 1286 => r := "10010100001101000010110101001000011";
      when 1287 => r := "10010100001101000010110010110100001";
      when 1288 => r := "10010100000101000010110000011111111";
      when 1289 => r := "10010100000101000010101110001011111";
      when 1290 => r := "10010100000001000010101011110111110";
      when 1291 => r := "10010100000001000010101001100011110";
      when 1292 => r := "10010011111001000010100111001111110";
      when 1293 => r := "10010011111001000010100100111011111";
      when 1294 => r := "10010011110001000010100010100111111";
      when 1295 => r := "10010011110001000010100000010100001";
      when 1296 => r := "10010011101001000010011110000000010";
      when 1297 => r := "10010011101001000010011011101100100";
      when 1298 => r := "10010011100101000010011001011001000";
      when 1299 => r := "10010011100101000010010111000101011";
      when 1300 => r := "10010011011101000010010100110001111";
      when 1301 => r := "10010011011101000010010010011110011";
      when 1302 => r := "10010011010101000010010000001011001";
      when 1303 => r := "10010011010101000010001101110111110";
      when 1304 => r := "10010011001101000010001011100100010";
      when 1305 => r := "10010011001101000010001001010001001";
      when 1306 => r := "10010011001001000010000110111101111";
      when 1307 => r := "10010011001001000010000100101010110";
      when 1308 => r := "10010011000001000010000010010111101";
      when 1309 => r := "10010011000001000010000000000100101";
      when 1310 => r := "10010010111001000001111101110001100";
      when 1311 => r := "10010010111001000001111011011110101";
      when 1312 => r := "10010010110001000001111001001011101";
      when 1313 => r := "10010010110001000001110110111000110";
      when 1314 => r := "10010010101101000001110100100110001";
      when 1315 => r := "10010010101101000001110010010011011";
      when 1316 => r := "10010010100101000001110000000000101";
      when 1317 => r := "10010010100101000001101101101110001";
      when 1318 => r := "10010010011101000001101011011011101";
      when 1319 => r := "10010010011101000001101001001001010";
      when 1320 => r := "10010010010101000001100110110110110";
      when 1321 => r := "10010010010101000001100100100100011";
      when 1322 => r := "10010010010001000001100010010001111";
      when 1323 => r := "10010010010001000001011111111111101";
      when 1324 => r := "10010010001001000001011101101101010";
      when 1325 => r := "10010010001001000001011011011011001";
      when 1326 => r := "10010010000001000001011001001001001";
      when 1327 => r := "10010010000001000001010110110111001";
      when 1328 => r := "10010001111001000001010100100101000";
      when 1329 => r := "10010001111001000001010010010011000";
      when 1330 => r := "10010001110101000001010000000001001";
      when 1331 => r := "10010001110101000001001101101111010";
      when 1332 => r := "10010001101101000001001011011101100";
      when 1333 => r := "10010001101101000001001001001011111";
      when 1334 => r := "10010001100101000001000110111010000";
      when 1335 => r := "10010001100101000001000100101000011";
      when 1336 => r := "10010001100001000001000010010110101";
      when 1337 => r := "10010001100001000001000000000101001";
      when 1338 => r := "10010001011001000000111101110011111";
      when 1339 => r := "10010001011001000000111011100010100";
      when 1340 => r := "10010001010001000000111001010001000";
      when 1341 => r := "10010001010001000000110110111111110";
      when 1342 => r := "10010001001001000000110100101110100";
      when 1343 => r := "10010001001001000000110010011101011";
      when 1344 => r := "10010001000101000000110000001100001";
      when 1345 => r := "10010001000101000000101101111011000";
      when 1346 => r := "10010000111101000000101011101001110";
      when 1347 => r := "10010000111101000000101001011000111";
      when 1348 => r := "10010000110101000000100111000111111";
      when 1349 => r := "10010000110101000000100100110111000";
      when 1350 => r := "10010000110001000000100010100110000";
      when 1351 => r := "10010000110001000000100000010101010";
      when 1352 => r := "10010000101001000000011110000100101";
      when 1353 => r := "10010000101001000000011011110100000";
      when 1354 => r := "10010000100001000000011001100011100";
      when 1355 => r := "10010000100001000000010111010010111";
      when 1356 => r := "10010000011101000000010101000010010";
      when 1357 => r := "10010000011101000000010010110001110";
      when 1358 => r := "10010000010101000000010000100001010";
      when 1359 => r := "10010000010101000000001110010001000";
      when 1360 => r := "10010000001101000000001100000000110";
      when 1361 => r := "10010000001101000000001001110000100";
      when 1362 => r := "10010000000101000000000111100000010";
      when 1363 => r := "10010000000101000000000101010000001";
      when 1364 => r := "10010000000001000000000011000000001";
      when 1365 => r := "10010000000001000000000000110000001";
      when 1366 => r := "10001111111000111111111110100000000";
      when 1367 => r := "10001111111000111111111100010000001";
      when 1368 => r := "10001111110000111111111010000000000";
      when 1369 => r := "10001111110000111111110111110000010";
      when 1370 => r := "10001111101100111111110101100000011";
      when 1371 => r := "10001111101100111111110011010000110";
      when 1372 => r := "10001111100100111111110001000001001";
      when 1373 => r := "10001111100100111111101110110001101";
      when 1374 => r := "10001111011100111111101100100010000";
      when 1375 => r := "10001111011100111111101010010010100";
      when 1376 => r := "10001111011000111111101000000010111";
      when 1377 => r := "10001111011000111111100101110011100";
      when 1378 => r := "10001111010000111111100011100100010";
      when 1379 => r := "10001111010000111111100001010101000";
      when 1380 => r := "10001111001000111111011111000101101";
      when 1381 => r := "10001111001000111111011100110110100";
      when 1382 => r := "10001111000100111111011010100111011";
      when 1383 => r := "10001111000100111111011000011000010";
      when 1384 => r := "10001110111100111111010110001001001";
      when 1385 => r := "10001110111100111111010011111010001";
      when 1386 => r := "10001110110100111111010001101011010";
      when 1387 => r := "10001110110100111111001111011100011";
      when 1388 => r := "10001110110000111111001101001101100";
      when 1389 => r := "10001110110000111111001010111110110";
      when 1390 => r := "10001110101000111111001000110000000";
      when 1391 => r := "10001110101000111111000110100001010";
      when 1392 => r := "10001110100000111111000100010010101";
      when 1393 => r := "10001110100000111111000010000100000";
      when 1394 => r := "10001110011100111110111111110101100";
      when 1395 => r := "10001110011100111110111101100111000";
      when 1396 => r := "10001110010100111110111011011000100";
      when 1397 => r := "10001110010100111110111001001010010";
      when 1398 => r := "10001110001100111110110110111100000";
      when 1399 => r := "10001110001100111110110100101101111";
      when 1400 => r := "10001110001000111110110010011111100";
      when 1401 => r := "10001110001000111110110000010001010";
      when 1402 => r := "10001110000000111110101110000011001";
      when 1403 => r := "10001110000000111110101011110101001";
      when 1404 => r := "10001101111000111110101001100111000";
      when 1405 => r := "10001101111000111110100111011001001";
      when 1406 => r := "10001101110100111110100101001011010";
      when 1407 => r := "10001101110100111110100010111101011";
      when 1408 => r := "10001101101100111110100000101111101";
      when 1409 => r := "10001101101100111110011110100001111";
      when 1410 => r := "10001101100100111110011100010100001";
      when 1411 => r := "10001101100100111110011010000110100";
      when 1412 => r := "10001101100000111110010111111001000";
      when 1413 => r := "10001101100000111110010101101011100";
      when 1414 => r := "10001101011000111110010011011101110";
      when 1415 => r := "10001101011000111110010001010000011";
      when 1416 => r := "10001101010100111110001111000010111";
      when 1417 => r := "10001101010100111110001100110101101";
      when 1418 => r := "10001101001100111110001010101000011";
      when 1419 => r := "10001101001100111110001000011011001";
      when 1420 => r := "10001101000100111110000110001110000";
      when 1421 => r := "10001101000100111110000100000000111";
      when 1422 => r := "10001101000000111110000001110011111";
      when 1423 => r := "10001101000000111101111111100110111";
      when 1424 => r := "10001100111000111101111101011001101";
      when 1425 => r := "10001100111000111101111011001100110";
      when 1426 => r := "10001100110000111101111001000000000";
      when 1427 => r := "10001100110000111101110110110011010";
      when 1428 => r := "10001100101100111101110100100110010";
      when 1429 => r := "10001100101100111101110010011001101";
      when 1430 => r := "10001100100100111101110000001101001";
      when 1431 => r := "10001100100100111101101110000000100";
      when 1432 => r := "10001100011100111101101011110011110";
      when 1433 => r := "10001100011100111101101001100111010";
      when 1434 => r := "10001100011000111101100111011010110";
      when 1435 => r := "10001100011000111101100101001110011";
      when 1436 => r := "10001100010000111101100011000001111";
      when 1437 => r := "10001100010000111101100000110101100";
      when 1438 => r := "10001100001100111101011110101001011";
      when 1439 => r := "10001100001100111101011100011101010";
      when 1440 => r := "10001100000100111101011010010001000";
      when 1441 => r := "10001100000100111101011000000100111";
      when 1442 => r := "10001011111100111101010101111000110";
      when 1443 => r := "10001011111100111101010011101100111";
      when 1444 => r := "10001011111000111101010001100000110";
      when 1445 => r := "10001011111000111101001111010100111";
      when 1446 => r := "10001011110000111101001101001001001";
      when 1447 => r := "10001011110000111101001010111101011";
      when 1448 => r := "10001011101000111101001000110001011";
      when 1449 => r := "10001011101000111101000110100101110";
      when 1450 => r := "10001011100100111101000100011010001";
      when 1451 => r := "10001011100100111101000010001110100";
      when 1452 => r := "10001011011100111101000000000010111";
      when 1453 => r := "10001011011100111100111101110111100";
      when 1454 => r := "10001011011000111100111011101100000";
      when 1455 => r := "10001011011000111100111001100000101";
      when 1456 => r := "10001011010000111100110111010101010";
      when 1457 => r := "10001011010000111100110101001010000";
      when 1458 => r := "10001011001000111100110010111110110";
      when 1459 => r := "10001011001000111100110000110011100";
      when 1460 => r := "10001011000100111100101110101000010";
      when 1461 => r := "10001011000100111100101100011101010";
      when 1462 => r := "10001010111100111100101010010010001";
      when 1463 => r := "10001010111100111100101000000111001";
      when 1464 => r := "10001010111000111100100101111100001";
      when 1465 => r := "10001010111000111100100011110001010";
      when 1466 => r := "10001010110000111100100001100110010";
      when 1467 => r := "10001010110000111100011111011011100";
      when 1468 => r := "10001010101000111100011101010000110";
      when 1469 => r := "10001010101000111100011011000110000";
      when 1470 => r := "10001010100100111100011000111011011";
      when 1471 => r := "10001010100100111100010110110000110";
      when 1472 => r := "10001010011100111100010100100110010";
      when 1473 => r := "10001010011100111100010010011011110";
      when 1474 => r := "10001010011000111100010000010001010";
      when 1475 => r := "10001010011000111100001110000110111";
      when 1476 => r := "10001010010000111100001011111100100";
      when 1477 => r := "10001010010000111100001001110010010";
      when 1478 => r := "10001010001100111100000111100111110";
      when 1479 => r := "10001010001100111100000101011101101";
      when 1480 => r := "10001010000100111100000011010011101";
      when 1481 => r := "10001010000100111100000001001001100";
      when 1482 => r := "10001001111100111011111110111111011";
      when 1483 => r := "10001001111100111011111100110101011";
      when 1484 => r := "10001001111000111011111010101011011";
      when 1485 => r := "10001001111000111011111000100001100";
      when 1486 => r := "10001001110000111011110110010111100";
      when 1487 => r := "10001001110000111011110100001101110";
      when 1488 => r := "10001001101100111011110010000100000";
      when 1489 => r := "10001001101100111011101111111010010";
      when 1490 => r := "10001001100100111011101101110000101";
      when 1491 => r := "10001001100100111011101011100111000";
      when 1492 => r := "10001001011100111011101001011101011";
      when 1493 => r := "10001001011100111011100111010011111";
      when 1494 => r := "10001001011000111011100101001010100";
      when 1495 => r := "10001001011000111011100011000001001";
      when 1496 => r := "10001001010000111011100000110111101";
      when 1497 => r := "10001001010000111011011110101110011";
      when 1498 => r := "10001001001100111011011100100101001";
      when 1499 => r := "10001001001100111011011010011011111";
      when 1500 => r := "10001001000100111011011000010010101";
      when 1501 => r := "10001001000100111011010110001001101";
      when 1502 => r := "10001001000000111011010100000000011";
      when 1503 => r := "10001001000000111011010001110111011";
      when 1504 => r := "10001000111000111011001111101110100";
      when 1505 => r := "10001000111000111011001101100101101";
      when 1506 => r := "10001000110000111011001011011100101";
      when 1507 => r := "10001000110000111011001001010011111";
      when 1508 => r := "10001000101100111011000111001011000";
      when 1509 => r := "10001000101100111011000101000010011";
      when 1510 => r := "10001000100100111011000010111001100";
      when 1511 => r := "10001000100100111011000000110001000";
      when 1512 => r := "10001000100000111010111110101000011";
      when 1513 => r := "10001000100000111010111100011111111";
      when 1514 => r := "10001000011000111010111010010111010";
      when 1515 => r := "10001000011000111010111000001110111";
      when 1516 => r := "10001000010100111010110110000110011";
      when 1517 => r := "10001000010100111010110011111110001";
      when 1518 => r := "10001000001100111010110001110101111";
      when 1519 => r := "10001000001100111010101111101101110";
      when 1520 => r := "10001000001000111010101101100101010";
      when 1521 => r := "10001000001000111010101011011101001";
      when 1522 => r := "10001000000000111010101001010101001";
      when 1523 => r := "10001000000000111010100111001101001";
      when 1524 => r := "10000111111000111010100101000101001";
      when 1525 => r := "10000111111000111010100010111101001";
      when 1526 => r := "10000111110100111010100000110101010";
      when 1527 => r := "10000111110100111010011110101101011";
      when 1528 => r := "10000111101100111010011100100101011";
      when 1529 => r := "10000111101100111010011010011101110";
      when 1530 => r := "10000111101000111010011000010101111";
      when 1531 => r := "10000111101000111010010110001110010";
      when 1532 => r := "10000111100000111010010100000110101";
      when 1533 => r := "10000111100000111010010001111111001";
      when 1534 => r := "10000111011100111010001111110111100";
      when 1535 => r := "10000111011100111010001101110000000";
      when 1536 => r := "10000111010100111010001011101000110";
      when 1537 => r := "10000111010100111010001001100001011";
      when 1538 => r := "10000111010000111010000111011010000";
      when 1539 => r := "10000111010000111010000101010010110";
      when 1540 => r := "10000111001000111010000011001011100";
      when 1541 => r := "10000111001000111010000001000100011";
      when 1542 => r := "10000111000100111001111110111101010";
      when 1543 => r := "10000111000100111001111100110110001";
      when 1544 => r := "10000110111100111001111010101111001";
      when 1545 => r := "10000110111100111001111000101000001";
      when 1546 => r := "10000110111000111001110110100001001";
      when 1547 => r := "10000110111000111001110100011010010";
      when 1548 => r := "10000110110000111001110010010011011";
      when 1549 => r := "10000110110000111001110000001100101";
      when 1550 => r := "10000110101000111001101110000101110";
      when 1551 => r := "10000110101000111001101011111111001";
      when 1552 => r := "10000110100100111001101001111000010";
      when 1553 => r := "10000110100100111001100111110001110";
      when 1554 => r := "10000110011100111001100101101011001";
      when 1555 => r := "10000110011100111001100011100100101";
      when 1556 => r := "10000110011000111001100001011110010";
      when 1557 => r := "10000110011000111001011111010111110";
      when 1558 => r := "10000110010000111001011101010001010";
      when 1559 => r := "10000110010000111001011011001011000";
      when 1560 => r := "10000110001100111001011001000100110";
      when 1561 => r := "10000110001100111001010110111110100";
      when 1562 => r := "10000110000100111001010100111000011";
      when 1563 => r := "10000110000100111001010010110010010";
      when 1564 => r := "10000110000000111001010000101100010";
      when 1565 => r := "10000110000000111001001110100110010";
      when 1566 => r := "10000101111000111001001100100000000";
      when 1567 => r := "10000101111000111001001010011010001";
      when 1568 => r := "10000101110100111001001000010100001";
      when 1569 => r := "10000101110100111001000110001110010";
      when 1570 => r := "10000101101100111001000100001000101";
      when 1571 => r := "10000101101100111001000010000010111";
      when 1572 => r := "10000101101000111000111111111101001";
      when 1573 => r := "10000101101000111000111101110111100";
      when 1574 => r := "10000101100000111000111011110001111";
      when 1575 => r := "10000101100000111000111001101100011";
      when 1576 => r := "10000101011100111000110111100110101";
      when 1577 => r := "10000101011100111000110101100001010";
      when 1578 => r := "10000101010100111000110011011100000";
      when 1579 => r := "10000101010100111000110001010110101";
      when 1580 => r := "10000101010000111000101111010001001";
      when 1581 => r := "10000101010000111000101101001011111";
      when 1582 => r := "10000101001000111000101011000110100";
      when 1583 => r := "10000101001000111000101001000001011";
      when 1584 => r := "10000101000100111000100110111100001";
      when 1585 => r := "10000101000100111000100100110111001";
      when 1586 => r := "10000100111100111000100010110010000";
      when 1587 => r := "10000100111100111000100000101101001";
      when 1588 => r := "10000100111000111000011110101000000";
      when 1589 => r := "10000100111000111000011100100011001";
      when 1590 => r := "10000100110000111000011010011110011";
      when 1591 => r := "10000100110000111000011000011001101";
      when 1592 => r := "10000100101100111000010110010100110";
      when 1593 => r := "10000100101100111000010100010000000";
      when 1594 => r := "10000100100100111000010010001011001";
      when 1595 => r := "10000100100100111000010000000110101";
      when 1596 => r := "10000100100000111000001110000010001";
      when 1597 => r := "10000100100000111000001011111101101";
      when 1598 => r := "10000100011000111000001001111001001";
      when 1599 => r := "10000100011000111000000111110100110";
      when 1600 => r := "10000100010100111000000101110000001";
      when 1601 => r := "10000100010100111000000011101011110";
      when 1602 => r := "10000100001100111000000001100111101";
      when 1603 => r := "10000100001100110111111111100011011";
      when 1604 => r := "10000100001000110111111101011111001";
      when 1605 => r := "10000100001000110111111011011011000";
      when 1606 => r := "10000100000000110111111001010110110";
      when 1607 => r := "10000100000000110111110111010010110";
      when 1608 => r := "10000011111100110111110101001110101";
      when 1609 => r := "10000011111100110111110011001010101";
      when 1610 => r := "10000011110100110111110001000110101";
      when 1611 => r := "10000011110100110111101111000010111";
      when 1612 => r := "10000011110000110111101100111110111";
      when 1613 => r := "10000011110000110111101010111011000";
      when 1614 => r := "10000011101000110111101000110111100";
      when 1615 => r := "10000011101000110111100110110011111";
      when 1616 => r := "10000011100100110111100100110000001";
      when 1617 => r := "10000011100100110111100010101100100";
      when 1618 => r := "10000011100000110111100000101000111";
      when 1619 => r := "10000011100000110111011110100101011";
      when 1620 => r := "10000011011000110111011100100001111";
      when 1621 => r := "10000011011000110111011010011110100";
      when 1622 => r := "10000011010100110111011000011011001";
      when 1623 => r := "10000011010100110111010110010111110";
      when 1624 => r := "10000011001100110111010100010100011";
      when 1625 => r := "10000011001100110111010010010001010";
      when 1626 => r := "10000011001000110111010000001101111";
      when 1627 => r := "10000011001000110111001110001010110";
      when 1628 => r := "10000011000000110111001100000111110";
      when 1629 => r := "10000011000000110111001010000100110";
      when 1630 => r := "10000010111100110111001000000001101";
      when 1631 => r := "10000010111100110111000101111110101";
      when 1632 => r := "10000010110100110111000011111011110";
      when 1633 => r := "10000010110100110111000001111001000";
      when 1634 => r := "10000010110000110110111111110101111";
      when 1635 => r := "10000010110000110110111101110011001";
      when 1636 => r := "10000010101000110110111011110000100";
      when 1637 => r := "10000010101000110110111001101101111";
      when 1638 => r := "10000010100100110110110111101011001";
      when 1639 => r := "10000010100100110110110101101000100";
      when 1640 => r := "10000010011100110110110011100101111";
      when 1641 => r := "10000010011100110110110001100011011";
      when 1642 => r := "10000010011000110110101111100001000";
      when 1643 => r := "10000010011000110110101101011110101";
      when 1644 => r := "10000010010000110110101011011100001";
      when 1645 => r := "10000010010000110110101001011001110";
      when 1646 => r := "10000010001100110110100111010111101";
      when 1647 => r := "10000010001100110110100101010101011";
      when 1648 => r := "10000010001000110110100011010011010";
      when 1649 => r := "10000010001000110110100001010001001";
      when 1650 => r := "10000010000000110110011111001110110";
      when 1651 => r := "10000010000000110110011101001100110";
      when 1652 => r := "10000001111100110110011011001010101";
      when 1653 => r := "10000001111100110110011001001000110";
      when 1654 => r := "10000001110100110110010111000110111";
      when 1655 => r := "10000001110100110110010101000101000";
      when 1656 => r := "10000001110000110110010011000011010";
      when 1657 => r := "10000001110000110110010001000001100";
      when 1658 => r := "10000001101000110110001110111111101";
      when 1659 => r := "10000001101000110110001100111101111";
      when 1660 => r := "10000001100100110110001010111100010";
      when 1661 => r := "10000001100100110110001000111010110";
      when 1662 => r := "10000001011100110110000110111001000";
      when 1663 => r := "10000001011100110110000100110111100";
      when 1664 => r := "10000001011000110110000010110110000";
      when 1665 => r := "10000001011000110110000000110100101";
      when 1666 => r := "10000001010100110101111110110011001";
      when 1667 => r := "10000001010100110101111100110001111";
      when 1668 => r := "10000001001100110101111010110000100";
      when 1669 => r := "10000001001100110101111000101111011";
      when 1670 => r := "10000001001000110101110110101110001";
      when 1671 => r := "10000001001000110101110100101101000";
      when 1672 => r := "10000001000000110101110010101011111";
      when 1673 => r := "10000001000000110101110000101010111";
      when 1674 => r := "10000000111100110101101110101001101";
      when 1675 => r := "10000000111100110101101100101000110";
      when 1676 => r := "10000000110100110101101010100111111";
      when 1677 => r := "10000000110100110101101000100111001";
      when 1678 => r := "10000000110000110101100110100110000";
      when 1679 => r := "10000000110000110101100100100101010";
      when 1680 => r := "10000000101100110101100010100100100";
      when 1681 => r := "10000000101100110101100000100011110";
      when 1682 => r := "10000000100100110101011110100011001";
      when 1683 => r := "10000000100100110101011100100010100";
      when 1684 => r := "10000000100000110101011010100010000";
      when 1685 => r := "10000000100000110101011000100001100";
      when 1686 => r := "10000000011000110101010110100000111";
      when 1687 => r := "10000000011000110101010100100000100";
      when 1688 => r := "10000000010100110101010010100000001";
      when 1689 => r := "10000000010100110101010000011111110";
      when 1690 => r := "10000000001100110101001110011111011";
      when 1691 => r := "10000000001100110101001100011111001";
      when 1692 => r := "10000000001000110101001010011111000";
      when 1693 => r := "10000000001000110101001000011110111";
      when 1694 => r := "10000000000100110101000110011110100";
      when 1695 => r := "10000000000100110101000100011110100";
      when 1696 => r := "01111111111100110101000010011110100";
      when 1697 => r := "01111111111100110101000000011110100";
      when 1698 => r := "01111111111000110100111110011110100";
      when 1699 => r := "01111111111000110100111100011110101";
      when 1700 => r := "01111111110000110100111010011110110";
      when 1701 => r := "01111111110000110100111000011111000";
      when 1702 => r := "01111111101100110100110110011111010";
      when 1703 => r := "01111111101100110100110100011111100";
      when 1704 => r := "01111111101000110100110010011111110";
      when 1705 => r := "01111111101000110100110000100000001";
      when 1706 => r := "01111111100000110100101110100000010";
      when 1707 => r := "01111111100000110100101100100000110";
      when 1708 => r := "01111111011100110100101010100001010";
      when 1709 => r := "01111111011100110100101000100001111";
      when 1710 => r := "01111111010100110100100110100010011";
      when 1711 => r := "01111111010100110100100100100011000";
      when 1712 => r := "01111111010000110100100010100011101";
      when 1713 => r := "01111111010000110100100000100100011";
      when 1714 => r := "01111111001100110100011110100101000";
      when 1715 => r := "01111111001100110100011100100101110";
      when 1716 => r := "01111111000100110100011010100110101";
      when 1717 => r := "01111111000100110100011000100111101";
      when 1718 => r := "01111111000000110100010110101000100";
      when 1719 => r := "01111111000000110100010100101001100";
      when 1720 => r := "01111110111000110100010010101010100";
      when 1721 => r := "01111110111000110100010000101011100";
      when 1722 => r := "01111110110100110100001110101100101";
      when 1723 => r := "01111110110100110100001100101101110";
      when 1724 => r := "01111110110000110100001010101110111";
      when 1725 => r := "01111110110000110100001000110000001";
      when 1726 => r := "01111110101000110100000110110001011";
      when 1727 => r := "01111110101000110100000100110010110";
      when 1728 => r := "01111110100100110100000010110100000";
      when 1729 => r := "01111110100100110100000000110101100";
      when 1730 => r := "01111110011100110011111110110111000";
      when 1731 => r := "01111110011100110011111100111000100";
      when 1732 => r := "01111110011000110011111010111001110";
      when 1733 => r := "01111110011000110011111000111011011";
      when 1734 => r := "01111110010100110011110110111101001";
      when 1735 => r := "01111110010100110011110100111110110";
      when 1736 => r := "01111110001100110011110011000000011";
      when 1737 => r := "01111110001100110011110001000010010";
      when 1738 => r := "01111110001000110011101111000100001";
      when 1739 => r := "01111110001000110011101101000110000";
      when 1740 => r := "01111110000000110011101011000111101";
      when 1741 => r := "01111110000000110011101001001001101";
      when 1742 => r := "01111101111100110011100111001011101";
      when 1743 => r := "01111101111100110011100101001101101";
      when 1744 => r := "01111101111000110011100011001111101";
      when 1745 => r := "01111101111000110011100001010001101";
      when 1746 => r := "01111101110000110011011111010011111";
      when 1747 => r := "01111101110000110011011101010110001";
      when 1748 => r := "01111101101100110011011011011000010";
      when 1749 => r := "01111101101100110011011001011010100";
      when 1750 => r := "01111101101000110011010111011100111";
      when 1751 => r := "01111101101000110011010101011111010";
      when 1752 => r := "01111101100000110011010011100001101";
      when 1753 => r := "01111101100000110011010001100100000";
      when 1754 => r := "01111101011100110011001111100110011";
      when 1755 => r := "01111101011100110011001101101000111";
      when 1756 => r := "01111101010100110011001011101011101";
      when 1757 => r := "01111101010100110011001001101110010";
      when 1758 => r := "01111101010000110011000111110000110";
      when 1759 => r := "01111101010000110011000101110011011";
      when 1760 => r := "01111101001100110011000011110110001";
      when 1761 => r := "01111101001100110011000001111000111";
      when 1762 => r := "01111101000100110010111111111011110";
      when 1763 => r := "01111101000100110010111101111110101";
      when 1764 => r := "01111101000000110010111100000001101";
      when 1765 => r := "01111101000000110010111010000100101";
      when 1766 => r := "01111100111100110010111000000111101";
      when 1767 => r := "01111100111100110010110110001010110";
      when 1768 => r := "01111100110100110010110100001101101";
      when 1769 => r := "01111100110100110010110010010000110";
      when 1770 => r := "01111100110000110010110000010011111";
      when 1771 => r := "01111100110000110010101110010111000";
      when 1772 => r := "01111100101100110010101100011010011";
      when 1773 => r := "01111100101100110010101010011101110";
      when 1774 => r := "01111100100100110010101000100000111";
      when 1775 => r := "01111100100100110010100110100100010";
      when 1776 => r := "01111100100000110010100100100111110";
      when 1777 => r := "01111100100000110010100010101011010";
      when 1778 => r := "01111100011000110010100000101110110";
      when 1779 => r := "01111100011000110010011110110010011";
      when 1780 => r := "01111100010100110010011100110101111";
      when 1781 => r := "01111100010100110010011010111001100";
      when 1782 => r := "01111100010000110010011000111101000";
      when 1783 => r := "01111100010000110010010111000000110";
      when 1784 => r := "01111100001000110010010101000100101";
      when 1785 => r := "01111100001000110010010011001000100";
      when 1786 => r := "01111100000100110010010001001100011";
      when 1787 => r := "01111100000100110010001111010000010";
      when 1788 => r := "01111100000000110010001101010100001";
      when 1789 => r := "01111100000000110010001011011000001";
      when 1790 => r := "01111011111000110010001001011100000";
      when 1791 => r := "01111011111000110010000111100000001";
      when 1792 => r := "01111011110100110010000101100100000";
      when 1793 => r := "01111011110100110010000011101000010";
      when 1794 => r := "01111011110000110010000001101100011";
      when 1795 => r := "01111011110000110001111111110000101";
      when 1796 => r := "01111011101000110001111101110101000";
      when 1797 => r := "01111011101000110001111011111001011";
      when 1798 => r := "01111011100100110001111001111101101";
      when 1799 => r := "01111011100100110001111000000010000";
      when 1800 => r := "01111011100000110001110110000110011";
      when 1801 => r := "01111011100000110001110100001010111";
      when 1802 => r := "01111011011000110001110010001111100";
      when 1803 => r := "01111011011000110001110000010100000";
      when 1804 => r := "01111011010100110001101110011000101";
      when 1805 => r := "01111011010100110001101100011101011";
      when 1806 => r := "01111011010000110001101010100001111";
      when 1807 => r := "01111011010000110001101000100110100";
      when 1808 => r := "01111011001000110001100110101011100";
      when 1809 => r := "01111011001000110001100100110000011";
      when 1810 => r := "01111011000100110001100010110101001";
      when 1811 => r := "01111011000100110001100000111010000";
      when 1812 => r := "01111011000000110001011110111110111";
      when 1813 => r := "01111011000000110001011101000011111";
      when 1814 => r := "01111010111000110001011011001000110";
      when 1815 => r := "01111010111000110001011001001101111";
      when 1816 => r := "01111010110100110001010111010011000";
      when 1817 => r := "01111010110100110001010101011000001";
      when 1818 => r := "01111010110000110001010011011101010";
      when 1819 => r := "01111010110000110001010001100010100";
      when 1820 => r := "01111010101000110001001111100111110";
      when 1821 => r := "01111010101000110001001101101101001";
      when 1822 => r := "01111010100100110001001011110010011";
      when 1823 => r := "01111010100100110001001001110111111";
      when 1824 => r := "01111010100000110001000111111101001";
      when 1825 => r := "01111010100000110001000110000010101";
      when 1826 => r := "01111010011000110001000100001000001";
      when 1827 => r := "01111010011000110001000010001101110";
      when 1828 => r := "01111010010100110001000000010011010";
      when 1829 => r := "01111010010100110000111110011000111";
      when 1830 => r := "01111010010000110000111100011110110";
      when 1831 => r := "01111010010000110000111010100100100";
      when 1832 => r := "01111010001000110000111000101010001";
      when 1833 => r := "01111010001000110000110110110000000";
      when 1834 => r := "01111010000100110000110100110101111";
      when 1835 => r := "01111010000100110000110010111011110";
      when 1836 => r := "01111010000000110000110001000001110";
      when 1837 => r := "01111010000000110000101111000111101";
      when 1838 => r := "01111001111000110000101101001101110";
      when 1839 => r := "01111001111000110000101011010011110";
      when 1840 => r := "01111001110100110000101001011001110";
      when 1841 => r := "01111001110100110000100111011111111";
      when 1842 => r := "01111001110000110000100101100110000";
      when 1843 => r := "01111001110000110000100011101100010";
      when 1844 => r := "01111001101000110000100001110010100";
      when 1845 => r := "01111001101000110000011111111000111";
      when 1846 => r := "01111001100100110000011101111111001";
      when 1847 => r := "01111001100100110000011100000101100";
      when 1848 => r := "01111001100000110000011010001100000";
      when 1849 => r := "01111001100000110000011000010010100";
      when 1850 => r := "01111001011100110000010110011000111";
      when 1851 => r := "01111001011100110000010100011111100";
      when 1852 => r := "01111001010100110000010010100110000";
      when 1853 => r := "01111001010100110000010000101100101";
      when 1854 => r := "01111001010000110000001110110011011";
      when 1855 => r := "01111001010000110000001100111010001";
      when 1856 => r := "01111001001100110000001011000000101";
      when 1857 => r := "01111001001100110000001001000111011";
      when 1858 => r := "01111001000100110000000111001110011";
      when 1859 => r := "01111001000100110000000101010101010";
      when 1860 => r := "01111001000000110000000011011100000";
      when 1861 => r := "01111001000000110000000001100011000";
      when 1862 => r := "01111000111100101111111111101010000";
      when 1863 => r := "01111000111100101111111101110001000";
      when 1864 => r := "01111000110100101111111011111000001";
      when 1865 => r := "01111000110100101111111001111111011";
      when 1866 => r := "01111000110000101111111000000110011";
      when 1867 => r := "01111000110000101111110110001101101";
      when 1868 => r := "01111000101100101111110100010100111";
      when 1869 => r := "01111000101100101111110010011100001";
      when 1870 => r := "01111000101000101111110000100011100";
      when 1871 => r := "01111000101000101111101110101010110";
      when 1872 => r := "01111000100000101111101100110010001";
      when 1873 => r := "01111000100000101111101010111001101";
      when 1874 => r := "01111000011100101111101001000001000";
      when 1875 => r := "01111000011100101111100111001000100";
      when 1876 => r := "01111000011000101111100101010000010";
      when 1877 => r := "01111000011000101111100011010111111";
      when 1878 => r := "01111000010000101111100001011111011";
      when 1879 => r := "01111000010000101111011111100111000";
      when 1880 => r := "01111000001100101111011101101110110";
      when 1881 => r := "01111000001100101111011011110110100";
      when 1882 => r := "01111000001000101111011001111110011";
      when 1883 => r := "01111000001000101111011000000110010";
      when 1884 => r := "01111000000100101111010110001110000";
      when 1885 => r := "01111000000100101111010100010101111";
      when 1886 => r := "01110111111100101111010010011101110";
      when 1887 => r := "01110111111100101111010000100101110";
      when 1888 => r := "01110111111000101111001110101101110";
      when 1889 => r := "01110111111000101111001100110101111";
      when 1890 => r := "01110111110100101111001010111110001";
      when 1891 => r := "01110111110100101111001001000110010";
      when 1892 => r := "01110111101100101111000111001110100";
      when 1893 => r := "01110111101100101111000101010110110";
      when 1894 => r := "01110111101000101111000011011111001";
      when 1895 => r := "01110111101000101111000001100111011";
      when 1896 => r := "01110111100100101110111111101111110";
      when 1897 => r := "01110111100100101110111101111000001";
      when 1898 => r := "01110111100000101110111100000000100";
      when 1899 => r := "01110111100000101110111010001001000";
      when 1900 => r := "01110111011000101110111000010001011";
      when 1901 => r := "01110111011000101110110110011010000";
      when 1902 => r := "01110111010100101110110100100010101";
      when 1903 => r := "01110111010100101110110010101011010";
      when 1904 => r := "01110111010000101110110000110011110";
      when 1905 => r := "01110111010000101110101110111100100";
      when 1906 => r := "01110111001000101110101101000101011";
      when 1907 => r := "01110111001000101110101011001110001";
      when 1908 => r := "01110111000100101110101001010110111";
      when 1909 => r := "01110111000100101110100111011111110";
      when 1910 => r := "01110111000000101110100101101000110";
      when 1911 => r := "01110111000000101110100011110001110";
      when 1912 => r := "01110110111100101110100001111010111";
      when 1913 => r := "01110110111100101110100000000011111";
      when 1914 => r := "01110110110100101110011110001100111";
      when 1915 => r := "01110110110100101110011100010110000";
      when 1916 => r := "01110110110000101110011010011111001";
      when 1917 => r := "01110110110000101110011000101000011";
      when 1918 => r := "01110110101100101110010110110001100";
      when 1919 => r := "01110110101100101110010100111010110";
      when 1920 => r := "01110110101000101110010011000100001";
      when 1921 => r := "01110110101000101110010001001101100";
      when 1922 => r := "01110110100000101110001111010110111";
      when 1923 => r := "01110110100000101110001101100000010";
      when 1924 => r := "01110110011100101110001011101001111";
      when 1925 => r := "01110110011100101110001001110011011";
      when 1926 => r := "01110110011000101110000111111100111";
      when 1927 => r := "01110110011000101110000110000110100";
      when 1928 => r := "01110110010100101110000100001111111";
      when 1929 => r := "01110110010100101110000010011001101";
      when 1930 => r := "01110110001100101110000000100011011";
      when 1931 => r := "01110110001100101101111110101101001";
      when 1932 => r := "01110110001000101101111100110111000";
      when 1933 => r := "01110110001000101101111011000000110";
      when 1934 => r := "01110110000100101101111001001010101";
      when 1935 => r := "01110110000100101101110111010100101";
      when 1936 => r := "01110110000000101101110101011110100";
      when 1937 => r := "01110110000000101101110011101000100";
      when 1938 => r := "01110101111000101101110001110010011";
      when 1939 => r := "01110101111000101101101111111100100";
      when 1940 => r := "01110101110100101101101110000110101";
      when 1941 => r := "01110101110100101101101100010000110";
      when 1942 => r := "01110101110000101101101010011011000";
      when 1943 => r := "01110101110000101101101000100101010";
      when 1944 => r := "01110101101100101101100110101111010";
      when 1945 => r := "01110101101100101101100100111001101";
      when 1946 => r := "01110101100100101101100011000100000";
      when 1947 => r := "01110101100100101101100001001110011";
      when 1948 => r := "01110101100000101101011111011000110";
      when 1949 => r := "01110101100000101101011101100011010";
      when 1950 => r := "01110101011100101101011011101101110";
      when 1951 => r := "01110101011100101101011001111000010";
      when 1952 => r := "01110101011000101101011000000010110";
      when 1953 => r := "01110101011000101101010110001101011";
      when 1954 => r := "01110101010000101101010100011000000";
      when 1955 => r := "01110101010000101101010010100010101";
      when 1956 => r := "01110101001100101101010000101101100";
      when 1957 => r := "01110101001100101101001110111000010";
      when 1958 => r := "01110101001000101101001101000010111";
      when 1959 => r := "01110101001000101101001011001101110";
      when 1960 => r := "01110101000100101101001001011000101";
      when 1961 => r := "01110101000100101101000111100011101";
      when 1962 => r := "01110100111100101101000101101110011";
      when 1963 => r := "01110100111100101101000011111001100";
      when 1964 => r := "01110100111000101101000010000100011";
      when 1965 => r := "01110100111000101101000000001111100";
      when 1966 => r := "01110100110100101100111110011010101";
      when 1967 => r := "01110100110100101100111100100101110";
      when 1968 => r := "01110100110000101100111010110001001";
      when 1969 => r := "01110100110000101100111000111100011";
      when 1970 => r := "01110100101000101100110111000111100";
      when 1971 => r := "01110100101000101100110101010010110";
      when 1972 => r := "01110100100100101100110011011110000";
      when 1973 => r := "01110100100100101100110001101001011";
      when 1974 => r := "01110100100000101100101111110101000";
      when 1975 => r := "01110100100000101100101110000000100";
      when 1976 => r := "01110100011100101100101100001011110";
      when 1977 => r := "01110100011100101100101010010111011";
      when 1978 => r := "01110100011000101100101000100010111";
      when 1979 => r := "01110100011000101100100110101110100";
      when 1980 => r := "01110100010000101100100100111010001";
      when 1981 => r := "01110100010000101100100011000101111";
      when 1982 => r := "01110100001100101100100001010001100";
      when 1983 => r := "01110100001100101100011111011101011";
      when 1984 => r := "01110100001000101100011101101001001";
      when 1985 => r := "01110100001000101100011011110101000";
      when 1986 => r := "01110100000100101100011010000000110";
      when 1987 => r := "01110100000100101100011000001100101";
      when 1988 => r := "01110011111100101100010110011000110";
      when 1989 => r := "01110011111100101100010100100100110";
      when 1990 => r := "01110011111000101100010010110000101";
      when 1991 => r := "01110011111000101100010000111100110";
      when 1992 => r := "01110011110100101100001111001000111";
      when 1993 => r := "01110011110100101100001101010101001";
      when 1994 => r := "01110011110000101100001011100001010";
      when 1995 => r := "01110011110000101100001001101101100";
      when 1996 => r := "01110011101100101100000111111001100";
      when 1997 => r := "01110011101100101100000110000101111";
      when 1998 => r := "01110011100100101100000100010010001";
      when 1999 => r := "01110011100100101100000010011110100";
      when 2000 => r := "01110011100000101100000000101011000";
      when 2001 => r := "01110011100000101011111110110111011";
      when 2002 => r := "01110011011100101011111101000011111";
      when 2003 => r := "01110011011100101011111011010000100";
      when 2004 => r := "01110011011000101011111001011101000";
      when 2005 => r := "01110011011000101011110111101001101";
      when 2006 => r := "01110011010000101011110101110110001";
      when 2007 => r := "01110011010000101011110100000010111";
      when 2008 => r := "01110011001100101011110010001111110";
      when 2009 => r := "01110011001100101011110000011100100";
      when 2010 => r := "01110011001000101011101110101001001";
      when 2011 => r := "01110011001000101011101100110110000";
      when 2012 => r := "01110011000100101011101011000010111";
      when 2013 => r := "01110011000100101011101001001111111";
      when 2014 => r := "01110011000000101011100111011100110";
      when 2015 => r := "01110011000000101011100101101001110";
      when 2016 => r := "01110010111000101011100011110110100";
      when 2017 => r := "01110010111000101011100010000011101";
      when 2018 => r := "01110010110100101011100000010000101";
      when 2019 => r := "01110010110100101011011110011101110";
      when 2020 => r := "01110010110000101011011100101011010";
      when 2021 => r := "01110010110000101011011010111000011";
      when 2022 => r := "01110010101100101011011001000101100";
      when 2023 => r := "01110010101100101011010111010010110";
      when 2024 => r := "01110010101000101011010101100000000";
      when 2025 => r := "01110010101000101011010011101101011";
      when 2026 => r := "01110010100000101011010001111010110";
      when 2027 => r := "01110010100000101011010000001000010";
      when 2028 => r := "01110010011100101011001110010101110";
      when 2029 => r := "01110010011100101011001100100011010";
      when 2030 => r := "01110010011000101011001010110000101";
      when 2031 => r := "01110010011000101011001000111110010";
      when 2032 => r := "01110010010100101011000111001011111";
      when 2033 => r := "01110010010100101011000101011001100";
      when 2034 => r := "01110010010000101011000011100111010";
      when 2035 => r := "01110010010000101011000001110101000";
      when 2036 => r := "01110010001000101011000000000010110";
      when 2037 => r := "01110010001000101010111110010000100";
      when 2038 => r := "01110010000100101010111100011110011";
      when 2039 => r := "01110010000100101010111010101100010";
      when 2040 => r := "01110010000000101010111000111010001";
      when 2041 => r := "01110010000000101010110111001000001";
      when 2042 => r := "01110001111100101010110101010110000";
      when 2043 => r := "01110001111100101010110011100100001";
      when 2044 => r := "01110001111000101010110001110010001";
      when 2045 => r := "01110001111000101010110000000000010";
      when 2046 => r := "01110001110100101010101110001110011";
      when 2047 => r := "01110001110100101010101100011100100";
      when 2048 => r := "01110001101100101010101010101010110";
      when 2049 => r := "01110001101100101010101000111001000";
      when 2050 => r := "01110001101000101010100111000111001";
      when 2051 => r := "01110001101000101010100101010101011";
      when 2052 => r := "01110001100100101010100011100011111";
      when 2053 => r := "01110001100100101010100001110010010";
      when 2054 => r := "01110001100000101010100000000000110";
      when 2055 => r := "01110001100000101010011110001111010";
      when 2056 => r := "01110001011100101010011100011101111";
      when 2057 => r := "01110001011100101010011010101100011";
      when 2058 => r := "01110001010100101010011000111010101";
      when 2059 => r := "01110001010100101010010111001001010";
      when 2060 => r := "01110001010000101010010101011000000";
      when 2061 => r := "01110001010000101010010011100110110";
      when 2062 => r := "01110001001100101010010001110101011";
      when 2063 => r := "01110001001100101010010000000100001";
      when 2064 => r := "01110001001000101010001110010010111";
      when 2065 => r := "01110001001000101010001100100001110";
      when 2066 => r := "01110001000100101010001010110000110";
      when 2067 => r := "01110001000100101010001000111111101";
      when 2068 => r := "01110001000000101010000111001110100";
      when 2069 => r := "01110001000000101010000101011101100";
      when 2070 => r := "01110000111000101010000011101100011";
      when 2071 => r := "01110000111000101010000001111011100";
      when 2072 => r := "01110000110100101010000000001010110";
      when 2073 => r := "01110000110100101001111110011001111";
      when 2074 => r := "01110000110000101001111100101001000";
      when 2075 => r := "01110000110000101001111010111000001";
      when 2076 => r := "01110000101100101001111001000111011";
      when 2077 => r := "01110000101100101001110111010110101";
      when 2078 => r := "01110000101000101001110101100101111";
      when 2079 => r := "01110000101000101001110011110101010";
      when 2080 => r := "01110000100100101001110010000100101";
      when 2081 => r := "01110000100100101001110000010100001";
      when 2082 => r := "01110000011100101001101110100011100";
      when 2083 => r := "01110000011100101001101100110011000";
      when 2084 => r := "01110000011000101001101011000010101";
      when 2085 => r := "01110000011000101001101001010010001";
      when 2086 => r := "01110000010100101001100111100001110";
      when 2087 => r := "01110000010100101001100101110001011";
      when 2088 => r := "01110000010000101001100100000001001";
      when 2089 => r := "01110000010000101001100010010000111";
      when 2090 => r := "01110000001100101001100000100000100";
      when 2091 => r := "01110000001100101001011110110000010";
      when 2092 => r := "01110000001000101001011101000000001";
      when 2093 => r := "01110000001000101001011011010000000";
      when 2094 => r := "01110000000000101001011001011111110";
      when 2095 => r := "01110000000000101001010111101111101";
      when 2096 => r := "01101111111100101001010101111111110";
      when 2097 => r := "01101111111100101001010100001111111";
      when 2098 => r := "01101111111000101001010010011111110";
      when 2099 => r := "01101111111000101001010000101111111";
      when 2100 => r := "01101111110100101001001110111111111";
      when 2101 => r := "01101111110100101001001101010000000";
      when 2102 => r := "01101111110000101001001011100000010";
      when 2103 => r := "01101111110000101001001001110000100";
      when 2104 => r := "01101111101100101001001000000000101";
      when 2105 => r := "01101111101100101001000110010001000";
      when 2106 => r := "01101111100100101001000100100001010";
      when 2107 => r := "01101111100100101001000010110001101";
      when 2108 => r := "01101111100000101001000001000010001";
      when 2109 => r := "01101111100000101000111111010010101";
      when 2110 => r := "01101111011100101000111101100010111";
      when 2111 => r := "01101111011100101000111011110011011";
      when 2112 => r := "01101111011000101000111010000011111";
      when 2113 => r := "01101111011000101000111000010100100";
      when 2114 => r := "01101111010100101000110110100101001";
      when 2115 => r := "01101111010100101000110100110101111";
      when 2116 => r := "01101111010000101000110011000110100";
      when 2117 => r := "01101111010000101000110001010111010";
      when 2118 => r := "01101111001100101000101111101000000";
      when 2119 => r := "01101111001100101000101101111000110";
      when 2120 => r := "01101111000100101000101100001001101";
      when 2121 => r := "01101111000100101000101010011010100";
      when 2122 => r := "01101111000000101000101000101011011";
      when 2123 => r := "01101111000000101000100110111100010";
      when 2124 => r := "01101110111100101000100101001101001";
      when 2125 => r := "01101110111100101000100011011110001";
      when 2126 => r := "01101110111000101000100001101111011";
      when 2127 => r := "01101110111000101000100000000000100";
      when 2128 => r := "01101110110100101000011110010001100";
      when 2129 => r := "01101110110100101000011100100010101";
      when 2130 => r := "01101110110000101000011010110011110";
      when 2131 => r := "01101110110000101000011001000101000";
      when 2132 => r := "01101110101100101000010111010110001";
      when 2133 => r := "01101110101100101000010101100111100";
      when 2134 => r := "01101110100100101000010011111001000";
      when 2135 => r := "01101110100100101000010010001010011";
      when 2136 => r := "01101110100000101000010000011011100";
      when 2137 => r := "01101110100000101000001110101101000";
      when 2138 => r := "01101110011100101000001100111110100";
      when 2139 => r := "01101110011100101000001011010000000";
      when 2140 => r := "01101110011000101000001001100001011";
      when 2141 => r := "01101110011000101000000111110011000";
      when 2142 => r := "01101110010100101000000110000100110";
      when 2143 => r := "01101110010100101000000100010110011";
      when 2144 => r := "01101110010000101000000010101000001";
      when 2145 => r := "01101110010000101000000000111001111";
      when 2146 => r := "01101110001100100111111111001011101";
      when 2147 => r := "01101110001100100111111101011101100";
      when 2148 => r := "01101110001000100111111011101111001";
      when 2149 => r := "01101110001000100111111010000001000";
      when 2150 => r := "01101110000000100111111000010010111";
      when 2151 => r := "01101110000000100111110110100100111";
      when 2152 => r := "01101101111100100111110100110110110";
      when 2153 => r := "01101101111100100111110011001000110";
      when 2154 => r := "01101101111000100111110001011010111";
      when 2155 => r := "01101101111000100111101111101100111";
      when 2156 => r := "01101101110100100111101101111111000";
      when 2157 => r := "01101101110100100111101100010001010";
      when 2158 => r := "01101101110000100111101010100011011";
      when 2159 => r := "01101101110000100111101000110101101";
      when 2160 => r := "01101101101100100111100111000111110";
      when 2161 => r := "01101101101100100111100101011010000";
      when 2162 => r := "01101101101000100111100011101100011";
      when 2163 => r := "01101101101000100111100001111110110";
      when 2164 => r := "01101101100100100111100000010001000";
      when 2165 => r := "01101101100100100111011110100011100";
      when 2166 => r := "01101101011100100111011100110101111";
      when 2167 => r := "01101101011100100111011011001000011";
      when 2168 => r := "01101101011000100111011001011010111";
      when 2169 => r := "01101101011000100111010111101101100";
      when 2170 => r := "01101101010100100111010110000000010";
      when 2171 => r := "01101101010100100111010100010010111";
      when 2172 => r := "01101101010000100111010010100101011";
      when 2173 => r := "01101101010000100111010000111000001";
      when 2174 => r := "01101101001100100111001111001010111";
      when 2175 => r := "01101101001100100111001101011101101";
      when 2176 => r := "01101101001000100111001011110000010";
      when 2177 => r := "01101101001000100111001010000011001";
      when 2178 => r := "01101101000100100111001000010110001";
      when 2179 => r := "01101101000100100111000110101001001";
      when 2180 => r := "01101101000000100111000100111011111";
      when 2181 => r := "01101101000000100111000011001110111";
      when 2182 => r := "01101100111100100111000001100010000";
      when 2183 => r := "01101100111100100110111111110101001";
      when 2184 => r := "01101100110100100110111110001000000";
      when 2185 => r := "01101100110100100110111100011011001";
      when 2186 => r := "01101100110000100110111010101110001";
      when 2187 => r := "01101100110000100110111001000001011";
      when 2188 => r := "01101100101100100110110111010100110";
      when 2189 => r := "01101100101100100110110101101000000";
      when 2190 => r := "01101100101000100110110011111011010";
      when 2191 => r := "01101100101000100110110010001110101";
      when 2192 => r := "01101100100100100110110000100001111";
      when 2193 => r := "01101100100100100110101110110101010";
      when 2194 => r := "01101100100000100110101101001000110";
      when 2195 => r := "01101100100000100110101011011100010";
      when 2196 => r := "01101100011100100110101001101111100";
      when 2197 => r := "01101100011100100110101000000011001";
      when 2198 => r := "01101100011000100110100110010110111";
      when 2199 => r := "01101100011000100110100100101010100";
      when 2200 => r := "01101100010100100110100010111110000";
      when 2201 => r := "01101100010100100110100001010001110";
      when 2202 => r := "01101100001100100110011111100101011";
      when 2203 => r := "01101100001100100110011101111001001";
      when 2204 => r := "01101100001000100110011100001100110";
      when 2205 => r := "01101100001000100110011010100000101";
      when 2206 => r := "01101100000100100110011000110100100";
      when 2207 => r := "01101100000100100110010111001000011";
      when 2208 => r := "01101100000000100110010101011100011";
      when 2209 => r := "01101100000000100110010011110000010";
      when 2210 => r := "01101011111100100110010010000100001";
      when 2211 => r := "01101011111100100110010000011000010";
      when 2212 => r := "01101011111000100110001110101100010";
      when 2213 => r := "01101011111000100110001101000000011";
      when 2214 => r := "01101011110100100110001011010100011";
      when 2215 => r := "01101011110100100110001001101000101";
      when 2216 => r := "01101011110000100110000111111100110";
      when 2217 => r := "01101011110000100110000110010001000";
      when 2218 => r := "01101011101100100110000100100101011";
      when 2219 => r := "01101011101100100110000010111001101";
      when 2220 => r := "01101011101000100110000001001110000";
      when 2221 => r := "01101011101000100101111111100010011";
      when 2222 => r := "01101011100100100101111101110110100";
      when 2223 => r := "01101011100100100101111100001010111";
      when 2224 => r := "01101011011100100101111010011111011";
      when 2225 => r := "01101011011100100101111000110011111";
      when 2226 => r := "01101011011000100101110111001000011";
      when 2227 => r := "01101011011000100101110101011101000";
      when 2228 => r := "01101011010100100101110011110001100";
      when 2229 => r := "01101011010100100101110010000110010";
      when 2230 => r := "01101011010000100101110000011010111";
      when 2231 => r := "01101011010000100101101110101111101";
      when 2232 => r := "01101011001100100101101101000100010";
      when 2233 => r := "01101011001100100101101011011001001";
      when 2234 => r := "01101011001000100101101001101101111";
      when 2235 => r := "01101011001000100101101000000010110";
      when 2236 => r := "01101011000100100101100110010111100";
      when 2237 => r := "01101011000100100101100100101100100";
      when 2238 => r := "01101011000000100101100011000001011";
      when 2239 => r := "01101011000000100101100001010110011";
      when 2240 => r := "01101010111100100101011111101011011";
      when 2241 => r := "01101010111100100101011110000000011";
      when 2242 => r := "01101010111000100101011100010101011";
      when 2243 => r := "01101010111000100101011010101010100";
      when 2244 => r := "01101010110100100101011000111111101";
      when 2245 => r := "01101010110100100101010111010100111";
      when 2246 => r := "01101010110000100101010101101010000";
      when 2247 => r := "01101010110000100101010011111111010";
      when 2248 => r := "01101010101000100101010010010100100";
      when 2249 => r := "01101010101000100101010000101001111";
      when 2250 => r := "01101010100100100101001110111111001";
      when 2251 => r := "01101010100100100101001101010100100";
      when 2252 => r := "01101010100000100101001011101001111";
      when 2253 => r := "01101010100000100101001001111111011";
      when 2254 => r := "01101010011100100101001000010100111";
      when 2255 => r := "01101010011100100101000110101010011";
      when 2256 => r := "01101010011000100101000100111111111";
      when 2257 => r := "01101010011000100101000011010101100";
      when 2258 => r := "01101010010100100101000001101011000";
      when 2259 => r := "01101010010100100101000000000000101";
      when 2260 => r := "01101010010000100100111110010110010";
      when 2261 => r := "01101010010000100100111100101100000";
      when 2262 => r := "01101010001100100100111011000001110";
      when 2263 => r := "01101010001100100100111001010111100";
      when 2264 => r := "01101010001000100100110111101101010";
      when 2265 => r := "01101010001000100100110110000011001";
      when 2266 => r := "01101010000100100100110100011001000";
      when 2267 => r := "01101010000100100100110010101111000";
      when 2268 => r := "01101010000000100100110001000100110";
      when 2269 => r := "01101010000000100100101111011010110";
      when 2270 => r := "01101001111100100100101101110000111";
      when 2271 => r := "01101001111100100100101100000110111";
      when 2272 => r := "01101001111000100100101010011100111";
      when 2273 => r := "01101001111000100100101000110011000";
      when 2274 => r := "01101001110100100100100111001001001";
      when 2275 => r := "01101001110100100100100101011111010";
      when 2276 => r := "01101001101100100100100011110101100";
      when 2277 => r := "01101001101100100100100010001011110";
      when 2278 => r := "01101001101000100100100000100010000";
      when 2279 => r := "01101001101000100100011110111000010";
      when 2280 => r := "01101001100100100100011101001110110";
      when 2281 => r := "01101001100100100100011011100101001";
      when 2282 => r := "01101001100000100100011001111011011";
      when 2283 => r := "01101001100000100100011000010001111";
      when 2284 => r := "01101001011100100100010110101000011";
      when 2285 => r := "01101001011100100100010100111110111";
      when 2286 => r := "01101001011000100100010011010101011";
      when 2287 => r := "01101001011000100100010001101011111";
      when 2288 => r := "01101001010100100100010000000010100";
      when 2289 => r := "01101001010100100100001110011001010";
      when 2290 => r := "01101001010000100100001100101111111";
      when 2291 => r := "01101001010000100100001011000110101";
      when 2292 => r := "01101001001100100100001001011101011";
      when 2293 => r := "01101001001100100100000111110100001";
      when 2294 => r := "01101001001000100100000110001010111";
      when 2295 => r := "01101001001000100100000100100001110";
      when 2296 => r := "01101001000100100100000010111000100";
      when 2297 => r := "01101001000100100100000001001111100";
      when 2298 => r := "01101001000000100011111111100110011";
      when 2299 => r := "01101001000000100011111101111101011";
      when 2300 => r := "01101000111100100011111100010100011";
      when 2301 => r := "01101000111100100011111010101011011";
      when 2302 => r := "01101000111000100011111001000010100";
      when 2303 => r := "01101000111000100011110111011001101";
      when 2304 => r := "01101000110100100011110101110000100";
      when 2305 => r := "01101000110100100011110100000111110";
      when 2306 => r := "01101000110000100011110010011110111";
      when 2307 => r := "01101000110000100011110000110110001";
      when 2308 => r := "01101000101100100011101111001101100";
      when 2309 => r := "01101000101100100011101101100100110";
      when 2310 => r := "01101000101000100011101011111100001";
      when 2311 => r := "01101000101000100011101010010011100";
      when 2312 => r := "01101000100100100011101000101011000";
      when 2313 => r := "01101000100100100011100111000010011";
      when 2314 => r := "01101000011100100011100101011001100";
      when 2315 => r := "01101000011100100011100011110001001";
      when 2316 => r := "01101000011000100011100010001000101";
      when 2317 => r := "01101000011000100011100000100000010";
      when 2318 => r := "01101000010100100011011110110111111";
      when 2319 => r := "01101000010100100011011101001111101";
      when 2320 => r := "01101000010000100011011011100111001";
      when 2321 => r := "01101000010000100011011001111110111";
      when 2322 => r := "01101000001100100011011000010110100";
      when 2323 => r := "01101000001100100011010110101110010";
      when 2324 => r := "01101000001000100011010101000110001";
      when 2325 => r := "01101000001000100011010011011110000";
      when 2326 => r := "01101000000100100011010001110101101";
      when 2327 => r := "01101000000100100011010000001101100";
      when 2328 => r := "01101000000000100011001110100101011";
      when 2329 => r := "01101000000000100011001100111101011";
      when 2330 => r := "01100111111100100011001011010101100";
      when 2331 => r := "01100111111100100011001001101101100";
      when 2332 => r := "01100111111000100011001000000101100";
      when 2333 => r := "01100111111000100011000110011101100";
      when 2334 => r := "01100111110100100011000100110101101";
      when 2335 => r := "01100111110100100011000011001101110";
      when 2336 => r := "01100111110000100011000001100101111";
      when 2337 => r := "01100111110000100010111111111110001";
      when 2338 => r := "01100111101100100010111110010110011";
      when 2339 => r := "01100111101100100010111100101110101";
      when 2340 => r := "01100111101000100010111011000111000";
      when 2341 => r := "01100111101000100010111001011111011";
      when 2342 => r := "01100111100100100010110111110111100";
      when 2343 => r := "01100111100100100010110110001111111";
      when 2344 => r := "01100111100000100010110100101000100";
      when 2345 => r := "01100111100000100010110011000000111";
      when 2346 => r := "01100111011100100010110001011001011";
      when 2347 => r := "01100111011100100010101111110001111";
      when 2348 => r := "01100111011000100010101110001010010";
      when 2349 => r := "01100111011000100010101100100010111";
      when 2350 => r := "01100111010100100010101010111011110";
      when 2351 => r := "01100111010100100010101001010100011";
      when 2352 => r := "01100111010000100010100111101101000";
      when 2353 => r := "01100111010000100010100110000101110";
      when 2354 => r := "01100111001100100010100100011110011";
      when 2355 => r := "01100111001100100010100010110111010";
      when 2356 => r := "01100111001000100010100001010000000";
      when 2357 => r := "01100111001000100010011111101000111";
      when 2358 => r := "01100111000100100010011110000001101";
      when 2359 => r := "01100111000100100010011100011010100";
      when 2360 => r := "01100111000000100010011010110011100";
      when 2361 => r := "01100111000000100010011001001100100";
      when 2362 => r := "01100110111100100010010111100101011";
      when 2363 => r := "01100110111100100010010101111110100";
      when 2364 => r := "01100110111000100010010100010111101";
      when 2365 => r := "01100110111000100010010010110000110";
      when 2366 => r := "01100110110100100010010001001001111";
      when 2367 => r := "01100110110100100010001111100011000";
      when 2368 => r := "01100110110000100010001101111100001";
      when 2369 => r := "01100110110000100010001100010101011";
      when 2370 => r := "01100110101100100010001010101110101";
      when 2371 => r := "01100110101100100010001001001000000";
      when 2372 => r := "01100110101000100010000111100001010";
      when 2373 => r := "01100110101000100010000101111010101";
      when 2374 => r := "01100110100100100010000100010100000";
      when 2375 => r := "01100110100100100010000010101101100";
      when 2376 => r := "01100110100000100010000001000111000";
      when 2377 => r := "01100110100000100001111111100000100";
      when 2378 => r := "01100110011100100001111101111001110";
      when 2379 => r := "01100110011100100001111100010011011";
      when 2380 => r := "01100110011000100001111010101101001";
      when 2381 => r := "01100110011000100001111001000110101";
      when 2382 => r := "01100110010100100001110111100000010";
      when 2383 => r := "01100110010100100001110101111010000";
      when 2384 => r := "01100110010000100001110100010011101";
      when 2385 => r := "01100110010000100001110010101101011";
      when 2386 => r := "01100110001100100001110001000111010";
      when 2387 => r := "01100110001100100001101111100001000";
      when 2388 => r := "01100110001000100001101101111010101";
      when 2389 => r := "01100110001000100001101100010100100";
      when 2390 => r := "01100110000100100001101010101110011";
      when 2391 => r := "01100110000100100001101001001000010";
      when 2392 => r := "01100110000000100001100111100010011";
      when 2393 => r := "01100110000000100001100101111100011";
      when 2394 => r := "01100101111100100001100100010110011";
      when 2395 => r := "01100101111100100001100010110000011";
      when 2396 => r := "01100101111000100001100001001010011";
      when 2397 => r := "01100101111000100001011111100100100";
      when 2398 => r := "01100101110100100001011101111110111";
      when 2399 => r := "01100101110100100001011100011001000";
      when 2400 => r := "01100101101100100001011010110011001";
      when 2401 => r := "01100101101100100001011001001101011";
      when 2402 => r := "01100101101000100001010111100111101";
      when 2403 => r := "01100101101000100001010110000001111";
      when 2404 => r := "01100101100100100001010100011100010";
      when 2405 => r := "01100101100100100001010010110110101";
      when 2406 => r := "01100101100000100001010001010001000";
      when 2407 => r := "01100101100000100001001111101011011";
      when 2408 => r := "01100101011100100001001110000101111";
      when 2409 => r := "01100101011100100001001100100000011";
      when 2410 => r := "01100101011000100001001010111010111";
      when 2411 => r := "01100101011000100001001001010101011";
      when 2412 => r := "01100101011000100001000111110000001";
      when 2413 => r := "01100101011000100001000110001010110";
      when 2414 => r := "01100101010100100001000100100101001";
      when 2415 => r := "01100101010100100001000010111111110";
      when 2416 => r := "01100101010000100001000001011010101";
      when 2417 => r := "01100101010000100000111111110101011";
      when 2418 => r := "01100101001100100000111110010000001";
      when 2419 => r := "01100101001100100000111100101010111";
      when 2420 => r := "01100101001000100000111011000101101";
      when 2421 => r := "01100101001000100000111001100000100";
      when 2422 => r := "01100101000100100000110111111011100";
      when 2423 => r := "01100101000100100000110110010110011";
      when 2424 => r := "01100101000000100000110100110001010";
      when 2425 => r := "01100101000000100000110011001100010";
      when 2426 => r := "01100100111100100000110001100111011";
      when 2427 => r := "01100100111100100000110000000010011";
      when 2428 => r := "01100100111000100000101110011101011";
      when 2429 => r := "01100100111000100000101100111000100";
      when 2430 => r := "01100100110100100000101011010011101";
      when 2431 => r := "01100100110100100000101001101110110";
      when 2432 => r := "01100100110000100000101000001010001";
      when 2433 => r := "01100100110000100000100110100101011";
      when 2434 => r := "01100100101100100000100101000000101";
      when 2435 => r := "01100100101100100000100011011100000";
      when 2436 => r := "01100100101000100000100001110111001";
      when 2437 => r := "01100100101000100000100000010010100";
      when 2438 => r := "01100100100100100000011110101101111";
      when 2439 => r := "01100100100100100000011101001001011";
      when 2440 => r := "01100100100000100000011011100100111";
      when 2441 => r := "01100100100000100000011010000000011";
      when 2442 => r := "01100100011100100000011000011011111";
      when 2443 => r := "01100100011100100000010110110111011";
      when 2444 => r := "01100100011000100000010101010011000";
      when 2445 => r := "01100100011000100000010011101110101";
      when 2446 => r := "01100100010100100000010010001010000";
      when 2447 => r := "01100100010100100000010000100101110";
      when 2448 => r := "01100100010000100000001111000001011";
      when 2449 => r := "01100100010000100000001101011101001";
      when 2450 => r := "01100100001100100000001011111001000";
      when 2451 => r := "01100100001100100000001010010100110";
      when 2452 => r := "01100100001000100000001000110000100";
      when 2453 => r := "01100100001000100000000111001100010";
      when 2454 => r := "01100100000100100000000101101000010";
      when 2455 => r := "01100100000100100000000100000100010";
      when 2456 => r := "01100100000000100000000010100000000";
      when 2457 => r := "01100100000000100000000000111100000";
      when 2458 => r := "01100011111100011111111111011000000";
      when 2459 => r := "01100011111100011111111101110100000";
      when 2460 => r := "01100011111000011111111100010000001";
      when 2461 => r := "01100011111000011111111010101100010";
      when 2462 => r := "01100011110100011111111001001000010";
      when 2463 => r := "01100011110100011111110111100100100";
      when 2464 => r := "01100011110000011111110110000000110";
      when 2465 => r := "01100011110000011111110100011101000";
      when 2466 => r := "01100011101100011111110010111001001";
      when 2467 => r := "01100011101100011111110001010101100";
      when 2468 => r := "01100011101000011111101111110001110";
      when 2469 => r := "01100011101000011111101110001110000";
      when 2470 => r := "01100011100100011111101100101010011";
      when 2471 => r := "01100011100100011111101011000110110";
      when 2472 => r := "01100011100000011111101001100011001";
      when 2473 => r := "01100011100000011111100111111111101";
      when 2474 => r := "01100011011100011111100110011100000";
      when 2475 => r := "01100011011100011111100100111000100";
      when 2476 => r := "01100011011000011111100011010101001";
      when 2477 => r := "01100011011000011111100001110001110";
      when 2478 => r := "01100011010100011111100000001110011";
      when 2479 => r := "01100011010100011111011110101011000";
      when 2480 => r := "01100011010000011111011101000111101";
      when 2481 => r := "01100011010000011111011011100100011";
      when 2482 => r := "01100011001100011111011010000000111";
      when 2483 => r := "01100011001100011111011000011101110";
      when 2484 => r := "01100011001000011111010110111010101";
      when 2485 => r := "01100011001000011111010101010111100";
      when 2486 => r := "01100011000100011111010011110100010";
      when 2487 => r := "01100011000100011111010010010001001";
      when 2488 => r := "01100011000000011111010000101110001";
      when 2489 => r := "01100011000000011111001111001011001";
      when 2490 => r := "01100010111100011111001101100111111";
      when 2491 => r := "01100010111100011111001100000101000";
      when 2492 => r := "01100010111000011111001010100010000";
      when 2493 => r := "01100010111000011111001000111111000";
      when 2494 => r := "01100010110100011111000111011100001";
      when 2495 => r := "01100010110100011111000101111001011";
      when 2496 => r := "01100010110000011111000100010110011";
      when 2497 => r := "01100010110000011111000010110011101";
      when 2498 => r := "01100010101100011111000001010000111";
      when 2499 => r := "01100010101100011110111111101110001";
      when 2500 => r := "01100010101100011110111110001011010";
      when 2501 => r := "01100010101100011110111100101000101";
      when 2502 => r := "01100010101000011110111011000101111";
      when 2503 => r := "01100010101000011110111001100011010";
      when 2504 => r := "01100010100100011110111000000000101";
      when 2505 => r := "01100010100100011110110110011110001";
      when 2506 => r := "01100010100000011110110100111011101";
      when 2507 => r := "01100010100000011110110011011001001";
      when 2508 => r := "01100010011100011110110001110110101";
      when 2509 => r := "01100010011100011110110000010100001";
      when 2510 => r := "01100010011000011110101110110001101";
      when 2511 => r := "01100010011000011110101101001111010";
      when 2512 => r := "01100010010100011110101011101100110";
      when 2513 => r := "01100010010100011110101010001010100";
      when 2514 => r := "01100010010000011110101000101000010";
      when 2515 => r := "01100010010000011110100111000110000";
      when 2516 => r := "01100010001100011110100101100011101";
      when 2517 => r := "01100010001100011110100100000001011";
      when 2518 => r := "01100010001000011110100010011111001";
      when 2519 => r := "01100010001000011110100000111101000";
      when 2520 => r := "01100010000100011110011111011010110";
      when 2521 => r := "01100010000100011110011101111000101";
      when 2522 => r := "01100010000000011110011100010110101";
      when 2523 => r := "01100010000000011110011010110100101";
      when 2524 => r := "01100001111100011110011001010010110";
      when 2525 => r := "01100001111100011110010111110000110";
      when 2526 => r := "01100001111000011110010110001110110";
      when 2527 => r := "01100001111000011110010100101100111";
      when 2528 => r := "01100001110100011110010011001010110";
      when 2529 => r := "01100001110100011110010001101000111";
      when 2530 => r := "01100001110000011110010000000111010";
      when 2531 => r := "01100001110000011110001110100101100";
      when 2532 => r := "01100001101100011110001101000011101";
      when 2533 => r := "01100001101100011110001011100001111";
      when 2534 => r := "01100001101000011110001010000000001";
      when 2535 => r := "01100001101000011110001000011110011";
      when 2536 => r := "01100001100100011110000110111100111";
      when 2537 => r := "01100001100100011110000101011011010";
      when 2538 => r := "01100001100000011110000011111001011";
      when 2539 => r := "01100001100000011110000010010111110";
      when 2540 => r := "01100001100000011110000000110110011";
      when 2541 => r := "01100001100000011101111111010100111";
      when 2542 => r := "01100001011100011101111101110011011";
      when 2543 => r := "01100001011100011101111100010001111";
      when 2544 => r := "01100001011000011101111010110000011";
      when 2545 => r := "01100001011000011101111001001111000";
      when 2546 => r := "01100001010100011101110111101101110";
      when 2547 => r := "01100001010100011101110110001100011";
      when 2548 => r := "01100001010000011101110100101011000";
      when 2549 => r := "01100001010000011101110011001001110";
      when 2550 => r := "01100001001100011101110001101000100";
      when 2551 => r := "01100001001100011101110000000111010";
      when 2552 => r := "01100001001000011101101110100110000";
      when 2553 => r := "01100001001000011101101101000100111";
      when 2554 => r := "01100001000100011101101011100011110";
      when 2555 => r := "01100001000100011101101010000010101";
      when 2556 => r := "01100001000000011101101000100001100";
      when 2557 => r := "01100001000000011101100111000000100";
      when 2558 => r := "01100000111100011101100101011111100";
      when 2559 => r := "01100000111100011101100011111110100";
      when 2560 => r := "01100000111000011101100010011101110";
      when 2561 => r := "01100000111000011101100000111100110";
      when 2562 => r := "01100000110100011101011111011011101";
      when 2563 => r := "01100000110100011101011101111010111";
      when 2564 => r := "01100000110000011101011100011010000";
      when 2565 => r := "01100000110000011101011010111001010";
      when 2566 => r := "01100000101100011101011001011000011";
      when 2567 => r := "01100000101100011101010111110111101";
      when 2568 => r := "01100000101000011101010110010110111";
      when 2569 => r := "01100000101000011101010100110110010";
      when 2570 => r := "01100000101000011101010011010101100";
      when 2571 => r := "01100000101000011101010001110100111";
      when 2572 => r := "01100000100100011101010000010100010";
      when 2573 => r := "01100000100100011101001110110011110";
      when 2574 => r := "01100000100000011101001101010011001";
      when 2575 => r := "01100000100000011101001011110010101";
      when 2576 => r := "01100000011100011101001010010010010";
      when 2577 => r := "01100000011100011101001000110001110";
      when 2578 => r := "01100000011000011101000111010001010";
      when 2579 => r := "01100000011000011101000101110000111";
      when 2580 => r := "01100000010100011101000100010000011";
      when 2581 => r := "01100000010100011101000010110000001";
      when 2582 => r := "01100000010000011101000001001111111";
      when 2583 => r := "01100000010000011100111111101111101";
      when 2584 => r := "01100000001100011100111110001111001";
      when 2585 => r := "01100000001100011100111100101111000";
      when 2586 => r := "01100000001000011100111011001110110";
      when 2587 => r := "01100000001000011100111001101110101";
      when 2588 => r := "01100000000100011100111000001110011";
      when 2589 => r := "01100000000100011100110110101110010";
      when 2590 => r := "01100000000000011100110101001110010";
      when 2591 => r := "01100000000000011100110011101110001";
      when 2592 => r := "01011111111100011100110010001110000";
      when 2593 => r := "01011111111100011100110000101110001";
      when 2594 => r := "01011111111000011100101111001110010";
      when 2595 => r := "01011111111000011100101101101110010";
      when 2596 => r := "01011111111000011100101100001110001";
      when 2597 => r := "01011111111000011100101010101110010";
      when 2598 => r := "01011111110100011100101001001110100";
      when 2599 => r := "01011111110100011100100111101110110";
      when 2600 => r := "01011111110000011100100110001110111";
      when 2601 => r := "01011111110000011100100100101111001";
      when 2602 => r := "01011111101100011100100011001111010";
      when 2603 => r := "01011111101100011100100001101111101";
      when 2604 => r := "01011111101000011100100000001111110";
      when 2605 => r := "01011111101000011100011110110000001";
      when 2606 => r := "01011111100100011100011101010000100";
      when 2607 => r := "01011111100100011100011011110000111";
      when 2608 => r := "01011111100000011100011010010001010";
      when 2609 => r := "01011111100000011100011000110001110";
      when 2610 => r := "01011111011100011100010111010010011";
      when 2611 => r := "01011111011100011100010101110010111";
      when 2612 => r := "01011111011000011100010100010011100";
      when 2613 => r := "01011111011000011100010010110100000";
      when 2614 => r := "01011111010100011100010001010100101";
      when 2615 => r := "01011111010100011100001111110101010";
      when 2616 => r := "01011111010000011100001110010110000";
      when 2617 => r := "01011111010000011100001100110110101";
      when 2618 => r := "01011111010000011100001011010111011";
      when 2619 => r := "01011111010000011100001001111000001";
      when 2620 => r := "01011111001100011100001000011000110";
      when 2621 => r := "01011111001100011100000110111001100";
      when 2622 => r := "01011111001000011100000101011010011";
      when 2623 => r := "01011111001000011100000011111011010";
      when 2624 => r := "01011111000100011100000010011100001";
      when 2625 => r := "01011111000100011100000000111101001";
      when 2626 => r := "01011111000000011011111111011101111";
      when 2627 => r := "01011111000000011011111101111110111";
      when 2628 => r := "01011110111100011011111100011111111";
      when 2629 => r := "01011110111100011011111011000001000";
      when 2630 => r := "01011110111000011011111001100001111";
      when 2631 => r := "01011110111000011011111000000010111";
      when 2632 => r := "01011110110100011011110110100100001";
      when 2633 => r := "01011110110100011011110101000101011";
      when 2634 => r := "01011110110000011011110011100110011";
      when 2635 => r := "01011110110000011011110010000111101";
      when 2636 => r := "01011110101100011011110000101000110";
      when 2637 => r := "01011110101100011011101111001010000";
      when 2638 => r := "01011110101000011011101101101011011";
      when 2639 => r := "01011110101000011011101100001100110";
      when 2640 => r := "01011110101000011011101010101110000";
      when 2641 => r := "01011110101000011011101001001111011";
      when 2642 => r := "01011110100100011011100111110000101";
      when 2643 => r := "01011110100100011011100110010010001";
      when 2644 => r := "01011110100000011011100100110011100";
      when 2645 => r := "01011110100000011011100011010101000";
      when 2646 => r := "01011110011100011011100001110110100";
      when 2647 => r := "01011110011100011011100000011000000";
      when 2648 => r := "01011110011000011011011110111001101";
      when 2649 => r := "01011110011000011011011101011011010";
      when 2650 => r := "01011110010100011011011011111100111";
      when 2651 => r := "01011110010100011011011010011110100";
      when 2652 => r := "01011110010000011011011001000000000";
      when 2653 => r := "01011110010000011011010111100001110";
      when 2654 => r := "01011110001100011011010110000011011";
      when 2655 => r := "01011110001100011011010100100101010";
      when 2656 => r := "01011110001000011011010011000111000";
      when 2657 => r := "01011110001000011011010001101000110";
      when 2658 => r := "01011110001000011011010000001010101";
      when 2659 => r := "01011110001000011011001110101100100";
      when 2660 => r := "01011110000100011011001101001110100";
      when 2661 => r := "01011110000100011011001011110000011";
      when 2662 => r := "01011110000000011011001010010010010";
      when 2663 => r := "01011110000000011011001000110100010";
      when 2664 => r := "01011101111100011011000111010110001";
      when 2665 => r := "01011101111100011011000101111000010";
      when 2666 => r := "01011101111000011011000100011010010";
      when 2667 => r := "01011101111000011011000010111100010";
      when 2668 => r := "01011101110100011011000001011110011";
      when 2669 => r := "01011101110100011011000000000000100";
      when 2670 => r := "01011101110000011010111110100010111";
      when 2671 => r := "01011101110000011010111101000101000";
      when 2672 => r := "01011101101100011010111011100111001";
      when 2673 => r := "01011101101100011010111010001001011";
      when 2674 => r := "01011101101000011010111000101011110";
      when 2675 => r := "01011101101000011010110111001110001";
      when 2676 => r := "01011101101000011010110101110000011";
      when 2677 => r := "01011101101000011010110100010010110";
      when 2678 => r := "01011101100100011010110010110101001";
      when 2679 => r := "01011101100100011010110001010111100";
      when 2680 => r := "01011101100000011010101111111010000";
      when 2681 => r := "01011101100000011010101110011100100";
      when 2682 => r := "01011101011100011010101100111110111";
      when 2683 => r := "01011101011100011010101011100001100";
      when 2684 => r := "01011101011000011010101010000100001";
      when 2685 => r := "01011101011000011010101000100110110";
      when 2686 => r := "01011101010100011010100111001001001";
      when 2687 => r := "01011101010100011010100101101011111";
      when 2688 => r := "01011101010000011010100100001110101";
      when 2689 => r := "01011101010000011010100010110001011";
      when 2690 => r := "01011101001100011010100001010100000";
      when 2691 => r := "01011101001100011010011111110110110";
      when 2692 => r := "01011101001000011010011110011001100";
      when 2693 => r := "01011101001000011010011100111100011";
      when 2694 => r := "01011101001000011010011011011111001";
      when 2695 => r := "01011101001000011010011010000010000";
      when 2696 => r := "01011101000100011010011000100100111";
      when 2697 => r := "01011101000100011010010111000111111";
      when 2698 => r := "01011101000000011010010101101010101";
      when 2699 => r := "01011101000000011010010100001101101";
      when 2700 => r := "01011100111100011010010010110000110";
      when 2701 => r := "01011100111100011010010001010011110";
      when 2702 => r := "01011100111000011010001111110110110";
      when 2703 => r := "01011100111000011010001110011001110";
      when 2704 => r := "01011100110100011010001100111100111";
      when 2705 => r := "01011100110100011010001011100000000";
      when 2706 => r := "01011100110000011010001010000011001";
      when 2707 => r := "01011100110000011010001000100110011";
      when 2708 => r := "01011100101100011010000111001001101";
      when 2709 => r := "01011100101100011010000101101100111";
      when 2710 => r := "01011100101100011010000100001111111";
      when 2711 => r := "01011100101100011010000010110011010";
      when 2712 => r := "01011100101000011010000001010110101";
      when 2713 => r := "01011100101000011001111111111010000";
      when 2714 => r := "01011100100100011001111110011101011";
      when 2715 => r := "01011100100100011001111101000000110";
      when 2716 => r := "01011100100000011001111011100100010";
      when 2717 => r := "01011100100000011001111010000111110";
      when 2718 => r := "01011100011100011001111000101011010";
      when 2719 => r := "01011100011100011001110111001110110";
      when 2720 => r := "01011100011000011001110101110010001";
      when 2721 => r := "01011100011000011001110100010101101";
      when 2722 => r := "01011100010100011001110010111001011";
      when 2723 => r := "01011100010100011001110001011101000";
      when 2724 => r := "01011100010100011001110000000000101";
      when 2725 => r := "01011100010100011001101110100100011";
      when 2726 => r := "01011100010000011001101101001000000";
      when 2727 => r := "01011100010000011001101011101011110";
      when 2728 => r := "01011100001100011001101010001111011";
      when 2729 => r := "01011100001100011001101000110011001";
      when 2730 => r := "01011100001000011001100111010111000";
      when 2731 => r := "01011100001000011001100101111010111";
      when 2732 => r := "01011100000100011001100100011110110";
      when 2733 => r := "01011100000100011001100011000010101";
      when 2734 => r := "01011100000000011001100001100110101";
      when 2735 => r := "01011100000000011001100000001010100";
      when 2736 => r := "01011011111100011001011110101110100";
      when 2737 => r := "01011011111100011001011101010010100";
      when 2738 => r := "01011011111000011001011011110110101";
      when 2739 => r := "01011011111000011001011010011010101";
      when 2740 => r := "01011011111000011001011000111110100";
      when 2741 => r := "01011011111000011001010111100010101";
      when 2742 => r := "01011011110100011001010110000110111";
      when 2743 => r := "01011011110100011001010100101011000";
      when 2744 => r := "01011011110000011001010011001111001";
      when 2745 => r := "01011011110000011001010001110011011";
      when 2746 => r := "01011011101100011001010000010111110";
      when 2747 => r := "01011011101100011001001110111100000";
      when 2748 => r := "01011011101000011001001101100000010";
      when 2749 => r := "01011011101000011001001100000100101";
      when 2750 => r := "01011011100100011001001010101000111";
      when 2751 => r := "01011011100100011001001001001101011";
      when 2752 => r := "01011011100000011001000111110001101";
      when 2753 => r := "01011011100000011001000110010110000";
      when 2754 => r := "01011011100000011001000100111010100";
      when 2755 => r := "01011011100000011001000011011111000";
      when 2756 => r := "01011011011100011001000010000011011";
      when 2757 => r := "01011011011100011001000000101000000";
      when 2758 => r := "01011011011000011000111111001100101";
      when 2759 => r := "01011011011000011000111101110001010";
      when 2760 => r := "01011011010100011000111100010101111";
      when 2761 => r := "01011011010100011000111010111010101";
      when 2762 => r := "01011011010000011000111001011111001";
      when 2763 => r := "01011011010000011000111000000011111";
      when 2764 => r := "01011011001100011000110110101000100";
      when 2765 => r := "01011011001100011000110101001101010";
      when 2766 => r := "01011011001000011000110011110010000";
      when 2767 => r := "01011011001000011000110010010110111";
      when 2768 => r := "01011011001000011000110000111011101";
      when 2769 => r := "01011011001000011000101111100000100";
      when 2770 => r := "01011011000100011000101110000101100";
      when 2771 => r := "01011011000100011000101100101010100";
      when 2772 => r := "01011011000000011000101011001111010";
      when 2773 => r := "01011011000000011000101001110100001";
      when 2774 => r := "01011010111100011000101000011001010";
      when 2775 => r := "01011010111100011000100110111110010";
      when 2776 => r := "01011010111000011000100101100011010";
      when 2777 => r := "01011010111000011000100100001000011";
      when 2778 => r := "01011010110100011000100010101101100";
      when 2779 => r := "01011010110100011000100001010010101";
      when 2780 => r := "01011010110100011000011111110111110";
      when 2781 => r := "01011010110100011000011110011100111";
      when 2782 => r := "01011010110000011000011101000010000";
      when 2783 => r := "01011010110000011000011011100111010";
      when 2784 => r := "01011010101100011000011010001100100";
      when 2785 => r := "01011010101100011000011000110001111";
      when 2786 => r := "01011010101000011000010111010111001";
      when 2787 => r := "01011010101000011000010101111100100";
      when 2788 => r := "01011010100100011000010100100001111";
      when 2789 => r := "01011010100100011000010011000111010";
      when 2790 => r := "01011010100000011000010001101100101";
      when 2791 => r := "01011010100000011000010000010010000";
      when 2792 => r := "01011010011100011000001110110111100";
      when 2793 => r := "01011010011100011000001101011101001";
      when 2794 => r := "01011010011100011000001100000010100";
      when 2795 => r := "01011010011100011000001010101000000";
      when 2796 => r := "01011010011000011000001001001101100";
      when 2797 => r := "01011010011000011000000111110011001";
      when 2798 => r := "01011010010100011000000110011000111";
      when 2799 => r := "01011010010100011000000100111110100";
      when 2800 => r := "01011010010000011000000011100100001";
      when 2801 => r := "01011010010000011000000010001001111";
      when 2802 => r := "01011010001100011000000000101111100";
      when 2803 => r := "01011010001100010111111111010101010";
      when 2804 => r := "01011010001000010111111101111011000";
      when 2805 => r := "01011010001000010111111100100000111";
      when 2806 => r := "01011010001000010111111011000110101";
      when 2807 => r := "01011010001000010111111001101100100";
      when 2808 => r := "01011010000100010111111000010010011";
      when 2809 => r := "01011010000100010111110110111000011";
      when 2810 => r := "01011010000000010111110101011110010";
      when 2811 => r := "01011010000000010111110100000100010";
      when 2812 => r := "01011001111100010111110010101010011";
      when 2813 => r := "01011001111100010111110001010000011";
      when 2814 => r := "01011001111000010111101111110110001";
      when 2815 => r := "01011001111000010111101110011100010";
      when 2816 => r := "01011001110100010111101101000010011";
      when 2817 => r := "01011001110100010111101011101000100";
      when 2818 => r := "01011001110100010111101010001110110";
      when 2819 => r := "01011001110100010111101000110100111";
      when 2820 => r := "01011001110000010111100111011011000";
      when 2821 => r := "01011001110000010111100110000001010";
      when 2822 => r := "01011001101100010111100100100111011";
      when 2823 => r := "01011001101100010111100011001101110";
      when 2824 => r := "01011001101000010111100001110100001";
      when 2825 => r := "01011001101000010111100000011010011";
      when 2826 => r := "01011001100100010111011111000000101";
      when 2827 => r := "01011001100100010111011101100111000";
      when 2828 => r := "01011001100000010111011100001101100";
      when 2829 => r := "01011001100000010111011010110100000";
      when 2830 => r := "01011001100000010111011001011010011";
      when 2831 => r := "01011001100000010111011000000000111";
      when 2832 => r := "01011001011100010111010110100111011";
      when 2833 => r := "01011001011100010111010101001110000";
      when 2834 => r := "01011001011000010111010011110100100";
      when 2835 => r := "01011001011000010111010010011011000";
      when 2836 => r := "01011001010100010111010001000001100";
      when 2837 => r := "01011001010100010111001111101000001";
      when 2838 => r := "01011001010000010111001110001111000";
      when 2839 => r := "01011001010000010111001100110101110";
      when 2840 => r := "01011001010000010111001011011100011";
      when 2841 => r := "01011001010000010111001010000011001";
      when 2842 => r := "01011001001100010111001000101001110";
      when 2843 => r := "01011001001100010111000111010000101";
      when 2844 => r := "01011001001000010111000101110111100";
      when 2845 => r := "01011001001000010111000100011110011";
      when 2846 => r := "01011001000100010111000011000101000";
      when 2847 => r := "01011001000100010111000001101100000";
      when 2848 => r := "01011001000000010111000000010011000";
      when 2849 => r := "01011001000000010110111110111010000";
      when 2850 => r := "01011000111100010110111101100000111";
      when 2851 => r := "01011000111100010110111100000111111";
      when 2852 => r := "01011000111100010110111010101110111";
      when 2853 => r := "01011000111100010110111001010110000";
      when 2854 => r := "01011000111000010110110111111101000";
      when 2855 => r := "01011000111000010110110110100100001";
      when 2856 => r := "01011000110100010110110101001011001";
      when 2857 => r := "01011000110100010110110011110010010";
      when 2858 => r := "01011000110000010110110010011001101";
      when 2859 => r := "01011000110000010110110001000000110";
      when 2860 => r := "01011000101100010110101111100111111";
      when 2861 => r := "01011000101100010110101110001111001";
      when 2862 => r := "01011000101100010110101100110110011";
      when 2863 => r := "01011000101100010110101011011101110";
      when 2864 => r := "01011000101000010110101010000101001";
      when 2865 => r := "01011000101000010110101000101100100";
      when 2866 => r := "01011000100100010110100111010011110";
      when 2867 => r := "01011000100100010110100101111011001";
      when 2868 => r := "01011000100000010110100100100010101";
      when 2869 => r := "01011000100000010110100011001010001";
      when 2870 => r := "01011000011100010110100001110001100";
      when 2871 => r := "01011000011100010110100000011001001";
      when 2872 => r := "01011000011000010110011111000000101";
      when 2873 => r := "01011000011000010110011101101000010";
      when 2874 => r := "01011000011000010110011100001111100";
      when 2875 => r := "01011000011000010110011010110111001";
      when 2876 => r := "01011000010100010110011001011110111";
      when 2877 => r := "01011000010100010110011000000110101";
      when 2878 => r := "01011000010000010110010110101110001";
      when 2879 => r := "01011000010000010110010101010101111";
      when 2880 => r := "01011000001100010110010011111101110";
      when 2881 => r := "01011000001100010110010010100101100";
      when 2882 => r := "01011000001000010110010001001101001";
      when 2883 => r := "01011000001000010110001111110100111";
      when 2884 => r := "01011000001000010110001110011100111";
      when 2885 => r := "01011000001000010110001101000100110";
      when 2886 => r := "01011000000100010110001011101100101";
      when 2887 => r := "01011000000100010110001010010100101";
      when 2888 => r := "01011000000000010110001000111100100";
      when 2889 => r := "01011000000000010110000111100100011";
      when 2890 => r := "01010111111100010110000110001100011";
      when 2891 => r := "01010111111100010110000100110100011";
      when 2892 => r := "01010111111000010110000011011100011";
      when 2893 => r := "01010111111000010110000010000100100";
      when 2894 => r := "01010111111000010110000000101100101";
      when 2895 => r := "01010111111000010101111111010100110";
      when 2896 => r := "01010111110100010101111101111100110";
      when 2897 => r := "01010111110100010101111100100101000";
      when 2898 => r := "01010111110000010101111011001101001";
      when 2899 => r := "01010111110000010101111001110101011";
      when 2900 => r := "01010111101100010101111000011101101";
      when 2901 => r := "01010111101100010101110111000101111";
      when 2902 => r := "01010111101000010101110101101110000";
      when 2903 => r := "01010111101000010101110100010110011";
      when 2904 => r := "01010111101000010101110010111110110";
      when 2905 => r := "01010111101000010101110001100111001";
      when 2906 => r := "01010111100100010101110000001111011";
      when 2907 => r := "01010111100100010101101110110111111";
      when 2908 => r := "01010111100000010101101101100000100";
      when 2909 => r := "01010111100000010101101100001001000";
      when 2910 => r := "01010111011100010101101010110001011";
      when 2911 => r := "01010111011100010101101001011010000";
      when 2912 => r := "01010111011000010101101000000010010";
      when 2913 => r := "01010111011000010101100110101010111";
      when 2914 => r := "01010111011000010101100101010011100";
      when 2915 => r := "01010111011000010101100011111100001";
      when 2916 => r := "01010111010100010101100010100100110";
      when 2917 => r := "01010111010100010101100001001101011";
      when 2918 => r := "01010111010000010101011111110110000";
      when 2919 => r := "01010111010000010101011110011110110";
      when 2920 => r := "01010111001100010101011101000111100";
      when 2921 => r := "01010111001100010101011011110000010";
      when 2922 => r := "01010111001000010101011010011001001";
      when 2923 => r := "01010111001000010101011001000001111";
      when 2924 => r := "01010111001000010101010111101010110";
      when 2925 => r := "01010111001000010101010110010011101";
      when 2926 => r := "01010111000100010101010100111100011";
      when 2927 => r := "01010111000100010101010011100101010";
      when 2928 => r := "01010111000000010101010010001110011";
      when 2929 => r := "01010111000000010101010000110111011";
      when 2930 => r := "01010110111100010101001111100000001";
      when 2931 => r := "01010110111100010101001110001001001";
      when 2932 => r := "01010110111000010101001100110010011";
      when 2933 => r := "01010110111000010101001011011011100";
      when 2934 => r := "01010110111000010101001010000100011";
      when 2935 => r := "01010110111000010101001000101101100";
      when 2936 => r := "01010110110100010101000111010110101";
      when 2937 => r := "01010110110100010101000101111111110";
      when 2938 => r := "01010110110000010101000100101001000";
      when 2939 => r := "01010110110000010101000011010010010";
      when 2940 => r := "01010110101100010101000001111011100";
      when 2941 => r := "01010110101100010101000000100100110";
      when 2942 => r := "01010110101000010100111111001110000";
      when 2943 => r := "01010110101000010100111101110111010";
      when 2944 => r := "01010110101000010100111100100000110";
      when 2945 => r := "01010110101000010100111011001010001";
      when 2946 => r := "01010110100100010100111001110011011";
      when 2947 => r := "01010110100100010100111000011100111";
      when 2948 => r := "01010110100000010100110111000110001";
      when 2949 => r := "01010110100000010100110101101111101";
      when 2950 => r := "01010110011100010100110100011001000";
      when 2951 => r := "01010110011100010100110011000010101";
      when 2952 => r := "01010110011100010100110001101100001";
      when 2953 => r := "01010110011100010100110000010101101";
      when 2954 => r := "01010110011000010100101110111111010";
      when 2955 => r := "01010110011000010100101101101000111";
      when 2956 => r := "01010110010100010100101100010010011";
      when 2957 => r := "01010110010100010100101010111100001";
      when 2958 => r := "01010110010000010100101001100101111";
      when 2959 => r := "01010110010000010100101000001111100";
      when 2960 => r := "01010110001100010100100110111001010";
      when 2961 => r := "01010110001100010100100101100011000";
      when 2962 => r := "01010110001100010100100100001100101";
      when 2963 => r := "01010110001100010100100010110110011";
      when 2964 => r := "01010110001000010100100001100000010";
      when 2965 => r := "01010110001000010100100000001010001";
      when 2966 => r := "01010110000100010100011110110100001";
      when 2967 => r := "01010110000100010100011101011110000";
      when 2968 => r := "01010110000000010100011100000111111";
      when 2969 => r := "01010110000000010100011010110001110";
      when 2970 => r := "01010101111100010100011001011011110";
      when 2971 => r := "01010101111100010100011000000101110";
      when 2972 => r := "01010101111100010100010110101111111";
      when 2973 => r := "01010101111100010100010101011001111";
      when 2974 => r := "01010101111000010100010100000011110";
      when 2975 => r := "01010101111000010100010010101101111";
      when 2976 => r := "01010101110100010100010001011000000";
      when 2977 => r := "01010101110100010100010000000010010";
      when 2978 => r := "01010101110000010100001110101100010";
      when 2979 => r := "01010101110000010100001101010110100";
      when 2980 => r := "01010101110000010100001100000000101";
      when 2981 => r := "01010101110000010100001010101010111";
      when 2982 => r := "01010101101100010100001001010101010";
      when 2983 => r := "01010101101100010100000111111111101";
      when 2984 => r := "01010101101000010100000110101001111";
      when 2985 => r := "01010101101000010100000101010100001";
      when 2986 => r := "01010101100100010100000011111110100";
      when 2987 => r := "01010101100100010100000010101000111";
      when 2988 => r := "01010101100000010100000001010011010";
      when 2989 => r := "01010101100000010011111111111101110";
      when 2990 => r := "01010101100000010011111110101000001";
      when 2991 => r := "01010101100000010011111101010010101";
      when 2992 => r := "01010101011100010011111011111101001";
      when 2993 => r := "01010101011100010011111010100111101";
      when 2994 => r := "01010101011000010011111001010010010";
      when 2995 => r := "01010101011000010011110111111100110";
      when 2996 => r := "01010101010100010011110110100111100";
      when 2997 => r := "01010101010100010011110101010010001";
      when 2998 => r := "01010101010100010011110011111100100";
      when 2999 => r := "01010101010100010011110010100111010";
      when 3000 => r := "01010101010000010011110001010010000";
      when 3001 => r := "01010101010000010011101111111100110";
      when 3002 => r := "01010101001100010011101110100111100";
      when 3003 => r := "01010101001100010011101101010010011";
      when 3004 => r := "01010101001000010011101011111101000";
      when 3005 => r := "01010101001000010011101010100111111";
      when 3006 => r := "01010101001000010011101001010010101";
      when 3007 => r := "01010101001000010011100111111101100";
      when 3008 => r := "01010101000100010011100110101000100";
      when 3009 => r := "01010101000100010011100101010011011";
      when 3010 => r := "01010101000000010011100011111110010";
      when 3011 => r := "01010101000000010011100010101001010";
      when 3012 => r := "01010100111100010011100001010100001";
      when 3013 => r := "01010100111100010011011111111111001";
      when 3014 => r := "01010100111000010011011110101010001";
      when 3015 => r := "01010100111000010011011101010101010";
      when 3016 => r := "01010100111000010011011100000000010";
      when 3017 => r := "01010100111000010011011010101011011";
      when 3018 => r := "01010100110100010011011001010110101";
      when 3019 => r := "01010100110100010011011000000001110";
      when 3020 => r := "01010100110000010011010110101100111";
      when 3021 => r := "01010100110000010011010101011000001";
      when 3022 => r := "01010100101100010011010100000011010";
      when 3023 => r := "01010100101100010011010010101110101";
      when 3024 => r := "01010100101100010011010001011001111";
      when 3025 => r := "01010100101100010011010000000101001";
      when 3026 => r := "01010100101000010011001110110000011";
      when 3027 => r := "01010100101000010011001101011011110";
      when 3028 => r := "01010100100100010011001100000111000";
      when 3029 => r := "01010100100100010011001010110010011";
      when 3030 => r := "01010100100000010011001001011101111";
      when 3031 => r := "01010100100000010011001000001001010";
      when 3032 => r := "01010100100000010011000110110100110";
      when 3033 => r := "01010100100000010011000101100000010";
      when 3034 => r := "01010100011100010011000100001011110";
      when 3035 => r := "01010100011100010011000010110111010";
      when 3036 => r := "01010100011000010011000001100010111";
      when 3037 => r := "01010100011000010011000000001110011";
      when 3038 => r := "01010100010100010010111110111001111";
      when 3039 => r := "01010100010100010010111101100101101";
      when 3040 => r := "01010100010100010010111100010001011";
      when 3041 => r := "01010100010100010010111010111101000";
      when 3042 => r := "01010100010000010010111001101000100";
      when 3043 => r := "01010100010000010010111000010100010";
      when 3044 => r := "01010100001100010010110111000000010";
      when 3045 => r := "01010100001100010010110101101100000";
      when 3046 => r := "01010100001000010010110100010111101";
      when 3047 => r := "01010100001000010010110011000011100";
      when 3048 => r := "01010100001000010010110001101111010";
      when 3049 => r := "01010100001000010010110000011011000";
      when 3050 => r := "01010100000100010010101111000111000";
      when 3051 => r := "01010100000100010010101101110010111";
      when 3052 => r := "01010100000000010010101100011110110";
      when 3053 => r := "01010100000000010010101011001010110";
      when 3054 => r := "01010011111100010010101001110110101";
      when 3055 => r := "01010011111100010010101000100010110";
      when 3056 => r := "01010011111100010010100111001110110";
      when 3057 => r := "01010011111100010010100101111010111";
      when 3058 => r := "01010011111000010010100100100110111";
      when 3059 => r := "01010011111000010010100011010011000";
      when 3060 => r := "01010011110100010010100001111111001";
      when 3061 => r := "01010011110100010010100000101011010";
      when 3062 => r := "01010011110000010010011111010111100";
      when 3063 => r := "01010011110000010010011110000011110";
      when 3064 => r := "01010011110000010010011100101111110";
      when 3065 => r := "01010011110000010010011011011100000";
      when 3066 => r := "01010011101100010010011010001000010";
      when 3067 => r := "01010011101100010010011000110100101";
      when 3068 => r := "01010011101000010010010111100000111";
      when 3069 => r := "01010011101000010010010110001101010";
      when 3070 => r := "01010011100100010010010100111001100";
      when 3071 => r := "01010011100100010010010011100101111";
      when 3072 => r := "01010011100100010010010010010010011";
      when 3073 => r := "01010011100100010010010000111110111";
      when 3074 => r := "01010011100000010010001111101011001";
      when 3075 => r := "01010011100000010010001110010111101";
      when 3076 => r := "01010011011100010010001101000100000";
      when 3077 => r := "01010011011100010010001011110000100";
      when 3078 => r := "01010011011000010010001010011101001";
      when 3079 => r := "01010011011000010010001001001001110";
      when 3080 => r := "01010011011000010010000111110110011";
      when 3081 => r := "01010011011000010010000110100011000";
      when 3082 => r := "01010011010100010010000101001111100";
      when 3083 => r := "01010011010100010010000011111100010";
      when 3084 => r := "01010011010000010010000010101000110";
      when 3085 => r := "01010011010000010010000001010101100";
      when 3086 => r := "01010011001100010010000000000010010";
      when 3087 => r := "01010011001100010001111110101111000";
      when 3088 => r := "01010011001100010001111101011011111";
      when 3089 => r := "01010011001100010001111100001000110";
      when 3090 => r := "01010011001000010001111010110101100";
      when 3091 => r := "01010011001000010001111001100010010";
      when 3092 => r := "01010011000100010001111000001111000";
      when 3093 => r := "01010011000100010001110110111011111";
      when 3094 => r := "01010011000000010001110101101000111";
      when 3095 => r := "01010011000000010001110100010101111";
      when 3096 => r := "01010011000000010001110011000010111";
      when 3097 => r := "01010011000000010001110001101111111";
      when 3098 => r := "01010010111100010001110000011100110";
      when 3099 => r := "01010010111100010001101111001001111";
      when 3100 => r := "01010010111000010001101101110110111";
      when 3101 => r := "01010010111000010001101100100011111";
      when 3102 => r := "01010010110100010001101011010001001";
      when 3103 => r := "01010010110100010001101001111110010";
      when 3104 => r := "01010010110100010001101000101011010";
      when 3105 => r := "01010010110100010001100111011000011";
      when 3106 => r := "01010010110000010001100110000101100";
      when 3107 => r := "01010010110000010001100100110010110";
      when 3108 => r := "01010010101100010001100011100000000";
      when 3109 => r := "01010010101100010001100010001101010";
      when 3110 => r := "01010010101100010001100000111010101";
      when 3111 => r := "01010010101100010001011111100111111";
      when 3112 => r := "01010010101000010001011110010101001";
      when 3113 => r := "01010010101000010001011101000010100";
      when 3114 => r := "01010010100100010001011011110000000";
      when 3115 => r := "01010010100100010001011010011101011";
      when 3116 => r := "01010010100000010001011001001010101";
      when 3117 => r := "01010010100000010001010111111000000";
      when 3118 => r := "01010010100000010001010110100101101";
      when 3119 => r := "01010010100000010001010101010011001";
      when 3120 => r := "01010010011100010001010100000000100";
      when 3121 => r := "01010010011100010001010010101110001";
      when 3122 => r := "01010010011000010001010001011011101";
      when 3123 => r := "01010010011000010001010000001001001";
      when 3124 => r := "01010010010100010001001110110110111";
      when 3125 => r := "01010010010100010001001101100100100";
      when 3126 => r := "01010010010100010001001100010010010";
      when 3127 => r := "01010010010100010001001010111111111";
      when 3128 => r := "01010010010000010001001001101101100";
      when 3129 => r := "01010010010000010001001000011011010";
      when 3130 => r := "01010010001100010001000111001001000";
      when 3131 => r := "01010010001100010001000101110110110";
      when 3132 => r := "01010010001000010001000100100100011";
      when 3133 => r := "01010010001000010001000011010010001";
      when 3134 => r := "01010010001000010001000010000000000";
      when 3135 => r := "01010010001000010001000000101101111";
      when 3136 => r := "01010010000100010000111111011011110";
      when 3137 => r := "01010010000100010000111110001001101";
      when 3138 => r := "01010010000000010000111100110111101";
      when 3139 => r := "01010010000000010000111011100101100";
      when 3140 => r := "01010010000000010000111010010011011";
      when 3141 => r := "01010010000000010000111001000001011";
      when 3142 => r := "01010001111100010000110111101111100";
      when 3143 => r := "01010001111100010000110110011101101";
      when 3144 => r := "01010001111000010000110101001011100";
      when 3145 => r := "01010001111000010000110011111001101";
      when 3146 => r := "01010001110100010000110010100111111";
      when 3147 => r := "01010001110100010000110001010110000";
      when 3148 => r := "01010001110100010000110000000100000";
      when 3149 => r := "01010001110100010000101110110010001";
      when 3150 => r := "01010001110000010000101101100000010";
      when 3151 => r := "01010001110000010000101100001110100";
      when 3152 => r := "01010001101100010000101010111100110";
      when 3153 => r := "01010001101100010000101001101011000";
      when 3154 => r := "01010001101100010000101000011001011";
      when 3155 => r := "01010001101100010000100111000111110";
      when 3156 => r := "01010001101000010000100101110101111";
      when 3157 => r := "01010001101000010000100100100100010";
      when 3158 => r := "01010001100100010000100011010010101";
      when 3159 => r := "01010001100100010000100010000001000";
      when 3160 => r := "01010001100000010000100000101111100";
      when 3161 => r := "01010001100000010000011111011101111";
      when 3162 => r := "01010001100000010000011110001100010";
      when 3163 => r := "01010001100000010000011100111010110";
      when 3164 => r := "01010001011100010000011011101001011";
      when 3165 => r := "01010001011100010000011010011000000";
      when 3166 => r := "01010001011000010000011001000110100";
      when 3167 => r := "01010001011000010000010111110101001";
      when 3168 => r := "01010001010100010000010110100011100";
      when 3169 => r := "01010001010100010000010101010010001";
      when 3170 => r := "01010001010100010000010100000000111";
      when 3171 => r := "01010001010100010000010010101111101";
      when 3172 => r := "01010001010000010000010001011110010";
      when 3173 => r := "01010001010000010000010000001100111";
      when 3174 => r := "01010001001100010000001110111011100";
      when 3175 => r := "01010001001100010000001101101010010";
      when 3176 => r := "01010001001100010000001100011001001";
      when 3177 => r := "01010001001100010000001011000111111";
      when 3178 => r := "01010001001000010000001001110110101";
      when 3179 => r := "01010001001000010000001000100101100";
      when 3180 => r := "01010001000100010000000111010100011";
      when 3181 => r := "01010001000100010000000110000011010";
      when 3182 => r := "01010001000000010000000100110010010";
      when 3183 => r := "01010001000000010000000011100001010";
      when 3184 => r := "01010001000000010000000010010000000";
      when 3185 => r := "01010001000000010000000000111111000";
      when 3186 => r := "01010000111100001111111111101110000";
      when 3187 => r := "01010000111100001111111110011101000";
      when 3188 => r := "01010000111000001111111101001100001";
      when 3189 => r := "01010000111000001111111011111011010";
      when 3190 => r := "01010000111000001111111010101010011";
      when 3191 => r := "01010000111000001111111001011001100";
      when 3192 => r := "01010000110100001111111000001000100";
      when 3193 => r := "01010000110100001111110110110111110";
      when 3194 => r := "01010000110000001111110101100110111";
      when 3195 => r := "01010000110000001111110100010110001";
      when 3196 => r := "01010000110000001111110011000101001";
      when 3197 => r := "01010000110000001111110001110100011";
      when 3198 => r := "01010000101100001111110000100011110";
      when 3199 => r := "01010000101100001111101111010011001";
      when 3200 => r := "01010000101000001111101110000010011";
      when 3201 => r := "01010000101000001111101100110001110";
      when 3202 => r := "01010000100100001111101011100000111";
      when 3203 => r := "01010000100100001111101010010000010";
      when 3204 => r := "01010000100100001111101000111111110";
      when 3205 => r := "01010000100100001111100111101111010";
      when 3206 => r := "01010000100000001111100110011110100";
      when 3207 => r := "01010000100000001111100101001110000";
      when 3208 => r := "01010000011100001111100011111101100";
      when 3209 => r := "01010000011100001111100010101101000";
      when 3210 => r := "01010000011100001111100001011100101";
      when 3211 => r := "01010000011100001111100000001100010";
      when 3212 => r := "01010000011000001111011110111011110";
      when 3213 => r := "01010000011000001111011101101011011";
      when 3214 => r := "01010000010100001111011100011010111";
      when 3215 => r := "01010000010100001111011011001010101";
      when 3216 => r := "01010000010000001111011001111010010";
      when 3217 => r := "01010000010000001111011000101010000";
      when 3218 => r := "01010000010000001111010111011001101";
      when 3219 => r := "01010000010000001111010110001001011";
      when 3220 => r := "01010000001100001111010100111001000";
      when 3221 => r := "01010000001100001111010011101000110";
      when 3222 => r := "01010000001000001111010010011000101";
      when 3223 => r := "01010000001000001111010001001000100";
      when 3224 => r := "01010000001000001111001111111000001";
      when 3225 => r := "01010000001000001111001110101000000";
      when 3226 => r := "01010000000100001111001101011000000";
      when 3227 => r := "01010000000100001111001100000111111";
      when 3228 => r := "01010000000000001111001010110111110";
      when 3229 => r := "01010000000000001111001001100111110";
      when 3230 => r := "01010000000000001111001000010111101";
      when 3231 => r := "01010000000000001111000111000111101";
      when 3232 => r := "01001111111100001111000101110111101";
      when 3233 => r := "01001111111100001111000100100111101";
      when 3234 => r := "01001111111000001111000011010111101";
      when 3235 => r := "01001111111000001111000010000111110";
      when 3236 => r := "01001111110100001111000000110111111";
      when 3237 => r := "01001111110100001110111111101000000";
      when 3238 => r := "01001111110100001110111110011000010";
      when 3239 => r := "01001111110100001110111101001000011";
      when 3240 => r := "01001111110000001110111011111000100";
      when 3241 => r := "01001111110000001110111010101000110";
      when 3242 => r := "01001111101100001110111001011001000";
      when 3243 => r := "01001111101100001110111000001001010";
      when 3244 => r := "01001111101100001110110110111001011";
      when 3245 => r := "01001111101100001110110101101001110";
      when 3246 => r := "01001111101000001110110100011001111";
      when 3247 => r := "01001111101000001110110011001010010";
      when 3248 => r := "01001111100100001110110001111010101";
      when 3249 => r := "01001111100100001110110000101011000";
      when 3250 => r := "01001111100100001110101111011011101";
      when 3251 => r := "01001111100100001110101110001100000";
      when 3252 => r := "01001111100000001110101100111100011";
      when 3253 => r := "01001111100000001110101011101100111";
      when 3254 => r := "01001111011100001110101010011101011";
      when 3255 => r := "01001111011100001110101001001101111";
      when 3256 => r := "01001111011100001110100111111110011";
      when 3257 => r := "01001111011100001110100110101110111";
      when 3258 => r := "01001111011000001110100101011111100";
      when 3259 => r := "01001111011000001110100100010000001";
      when 3260 => r := "01001111010100001110100011000000101";
      when 3261 => r := "01001111010100001110100001110001010";
      when 3262 => r := "01001111010000001110100000100010000";
      when 3263 => r := "01001111010000001110011111010010101";
      when 3264 => r := "01001111010000001110011110000011100";
      when 3265 => r := "01001111010000001110011100110100010";
      when 3266 => r := "01001111001100001110011011100100111";
      when 3267 => r := "01001111001100001110011010010101101";
      when 3268 => r := "01001111001000001110011001000110011";
      when 3269 => r := "01001111001000001110010111110111010";
      when 3270 => r := "01001111001000001110010110101000000";
      when 3271 => r := "01001111001000001110010101011000111";
      when 3272 => r := "01001111000100001110010100001001110";
      when 3273 => r := "01001111000100001110010010111010101";
      when 3274 => r := "01001111000000001110010001101011100";
      when 3275 => r := "01001111000000001110010000011100011";
      when 3276 => r := "01001111000000001110001111001101100";
      when 3277 => r := "01001111000000001110001101111110100";
      when 3278 => r := "01001110111100001110001100101111011";
      when 3279 => r := "01001110111100001110001011100000100";
      when 3280 => r := "01001110111000001110001010010001100";
      when 3281 => r := "01001110111000001110001001000010101";
      when 3282 => r := "01001110111000001110000111110011101";
      when 3283 => r := "01001110111000001110000110100100110";
      when 3284 => r := "01001110110100001110000101010101111";
      when 3285 => r := "01001110110100001110000100000111000";
      when 3286 => r := "01001110110000001110000010111000001";
      when 3287 => r := "01001110110000001110000001101001011";
      when 3288 => r := "01001110110000001110000000011010101";
      when 3289 => r := "01001110110000001101111111001011111";
      when 3290 => r := "01001110101100001101111101111101010";
      when 3291 => r := "01001110101100001101111100101110100";
      when 3292 => r := "01001110101000001101111011011111110";
      when 3293 => r := "01001110101000001101111010010001001";
      when 3294 => r := "01001110100100001101111001000010100";
      when 3295 => r := "01001110100100001101110111110100000";
      when 3296 => r := "01001110100100001101110110100101010";
      when 3297 => r := "01001110100100001101110101010110101";
      when 3298 => r := "01001110100000001101110100000111111";
      when 3299 => r := "01001110100000001101110010111001011";
      when 3300 => r := "01001110011100001101110001101010111";
      when 3301 => r := "01001110011100001101110000011100011";
      when 3302 => r := "01001110011100001101101111001110000";
      when 3303 => r := "01001110011100001101101101111111100";
      when 3304 => r := "01001110011000001101101100110001000";
      when 3305 => r := "01001110011000001101101011100010100";
      when 3306 => r := "01001110010100001101101010010100010";
      when 3307 => r := "01001110010100001101101001000101111";
      when 3308 => r := "01001110010100001101100111110111011";
      when 3309 => r := "01001110010100001101100110101001001";
      when 3310 => r := "01001110010000001101100101011010111";
      when 3311 => r := "01001110010000001101100100001100100";
      when 3312 => r := "01001110001100001101100010111110010";
      when 3313 => r := "01001110001100001101100001110000001";
      when 3314 => r := "01001110001100001101100000100001110";
      when 3315 => r := "01001110001100001101011111010011100";
      when 3316 => r := "01001110001000001101011110000101011";
      when 3317 => r := "01001110001000001101011100110111010";
      when 3318 => r := "01001110000100001101011011101001000";
      when 3319 => r := "01001110000100001101011010011010111";
      when 3320 => r := "01001110000100001101011001001100101";
      when 3321 => r := "01001110000100001101010111111110101";
      when 3322 => r := "01001110000000001101010110110000110";
      when 3323 => r := "01001110000000001101010101100010110";
      when 3324 => r := "01001101111100001101010100010100101";
      when 3325 => r := "01001101111100001101010011000110101";
      when 3326 => r := "01001101111100001101010001111000110";
      when 3327 => r := "01001101111100001101010000101010110";
      when 3328 => r := "01001101111000001101001111011100101";
      when 3329 => r := "01001101111000001101001110001110110";
      when 3330 => r := "01001101110100001101001101000000111";
      when 3331 => r := "01001101110100001101001011110011000";
      when 3332 => r := "01001101110100001101001010100101001";
      when 3333 => r := "01001101110100001101001001010111011";
      when 3334 => r := "01001101110000001101001000001001100";
      when 3335 => r := "01001101110000001101000110111011110";
      when 3336 => r := "01001101101100001101000101101110000";
      when 3337 => r := "01001101101100001101000100100000011";
      when 3338 => r := "01001101101100001101000011010010100";
      when 3339 => r := "01001101101100001101000010000100110";
      when 3340 => r := "01001101101000001101000000110111001";
      when 3341 => r := "01001101101000001100111111101001100";
      when 3342 => r := "01001101100100001100111110011011111";
      when 3343 => r := "01001101100100001100111101001110010";
      when 3344 => r := "01001101100100001100111100000000101";
      when 3345 => r := "01001101100100001100111010110011001";
      when 3346 => r := "01001101100000001100111001100101011";
      when 3347 => r := "01001101100000001100111000010111111";
      when 3348 => r := "01001101011100001100110111001010010";
      when 3349 => r := "01001101011100001100110101111100110";
      when 3350 => r := "01001101011100001100110100101111011";
      when 3351 => r := "01001101011100001100110011100001111";
      when 3352 => r := "01001101011000001100110010010100101";
      when 3353 => r := "01001101011000001100110001000111010";
      when 3354 => r := "01001101010100001100101111111001110";
      when 3355 => r := "01001101010100001100101110101100011";
      when 3356 => r := "01001101010100001100101101011111000";
      when 3357 => r := "01001101010100001100101100010001101";
      when 3358 => r := "01001101010000001100101011000100010";
      when 3359 => r := "01001101010000001100101001110111000";
      when 3360 => r := "01001101001100001100101000101001111";
      when 3361 => r := "01001101001100001100100111011100101";
      when 3362 => r := "01001101001100001100100110001111011";
      when 3363 => r := "01001101001100001100100101000010010";
      when 3364 => r := "01001101001000001100100011110100111";
      when 3365 => r := "01001101001000001100100010100111110";
      when 3366 => r := "01001101000100001100100001011010101";
      when 3367 => r := "01001101000100001100100000001101100";
      when 3368 => r := "01001101000100001100011111000000011";
      when 3369 => r := "01001101000100001100011101110011010";
      when 3370 => r := "01001101000000001100011100100110010";
      when 3371 => r := "01001101000000001100011011011001010";
      when 3372 => r := "01001100111100001100011010001100001";
      when 3373 => r := "01001100111100001100011000111111001";
      when 3374 => r := "01001100111100001100010111110010001";
      when 3375 => r := "01001100111100001100010110100101001";
      when 3376 => r := "01001100111000001100010101011000010";
      when 3377 => r := "01001100111000001100010100001011010";
      when 3378 => r := "01001100110100001100010010111110101";
      when 3379 => r := "01001100110100001100010001110001110";
      when 3380 => r := "01001100110100001100010000100100111";
      when 3381 => r := "01001100110100001100001111011000000";
      when 3382 => r := "01001100110000001100001110001011001";
      when 3383 => r := "01001100110000001100001100111110010";
      when 3384 => r := "01001100101100001100001011110001011";
      when 3385 => r := "01001100101100001100001010100100101";
      when 3386 => r := "01001100101100001100001001010111111";
      when 3387 => r := "01001100101100001100001000001011010";
      when 3388 => r := "01001100101000001100000110111110101";
      when 3389 => r := "01001100101000001100000101110010000";
      when 3390 => r := "01001100100100001100000100100101010";
      when 3391 => r := "01001100100100001100000011011000101";
      when 3392 => r := "01001100100100001100000010001100000";
      when 3393 => r := "01001100100100001100000000111111100";
      when 3394 => r := "01001100100000001011111111110011000";
      when 3395 => r := "01001100100000001011111110100110011";
      when 3396 => r := "01001100011100001011111101011001111";
      when 3397 => r := "01001100011100001011111100001101011";
      when 3398 => r := "01001100011100001011111011000000111";
      when 3399 => r := "01001100011100001011111001110100011";
      when 3400 => r := "01001100011000001011111000100111111";
      when 3401 => r := "01001100011000001011110111011011011";
      when 3402 => r := "01001100011000001011110110001111000";
      when 3403 => r := "01001100011000001011110101000010101";
      when 3404 => r := "01001100010100001011110011110110010";
      when 3405 => r := "01001100010100001011110010101010000";
      when 3406 => r := "01001100010000001011110001011101110";
      when 3407 => r := "01001100010000001011110000010001011";
      when 3408 => r := "01001100010000001011101111000101001";
      when 3409 => r := "01001100010000001011101101111000111";
      when 3410 => r := "01001100001100001011101100101100101";
      when 3411 => r := "01001100001100001011101011100000100";
      when 3412 => r := "01001100001000001011101010010100001";
      when 3413 => r := "01001100001000001011101001001000000";
      when 3414 => r := "01001100001000001011100111111011110";
      when 3415 => r := "01001100001000001011100110101111101";
      when 3416 => r := "01001100000100001011100101100011100";
      when 3417 => r := "01001100000100001011100100010111011";
      when 3418 => r := "01001100000000001011100011001011011";
      when 3419 => r := "01001100000000001011100001111111011";
      when 3420 => r := "01001100000000001011100000110011010";
      when 3421 => r := "01001100000000001011011111100111010";
      when 3422 => r := "01001011111100001011011110011011010";
      when 3423 => r := "01001011111100001011011101001111010";
      when 3424 => r := "01001011111000001011011100000011010";
      when 3425 => r := "01001011111000001011011010110111011";
      when 3426 => r := "01001011111000001011011001101011011";
      when 3427 => r := "01001011111000001011011000011111100";
      when 3428 => r := "01001011110100001011010111010011101";
      when 3429 => r := "01001011110100001011010110000111110";
      when 3430 => r := "01001011110000001011010100111011111";
      when 3431 => r := "01001011110000001011010011110000000";
      when 3432 => r := "01001011110000001011010010100100011";
      when 3433 => r := "01001011110000001011010001011000101";
      when 3434 => r := "01001011101100001011010000001100101";
      when 3435 => r := "01001011101100001011001111000001000";
      when 3436 => r := "01001011101000001011001101110101100";
      when 3437 => r := "01001011101000001011001100101001110";
      when 3438 => r := "01001011101000001011001011011110000";
      when 3439 => r := "01001011101000001011001010010010011";
      when 3440 => r := "01001011100100001011001001000110101";
      when 3441 => r := "01001011100100001011000111111011000";
      when 3442 => r := "01001011100100001011000110101111100";
      when 3443 => r := "01001011100100001011000101100011111";
      when 3444 => r := "01001011100000001011000100011000011";
      when 3445 => r := "01001011100000001011000011001100111";
      when 3446 => r := "01001011011100001011000010000001010";
      when 3447 => r := "01001011011100001011000000110101110";
      when 3448 => r := "01001011011100001010111111101010011";
      when 3449 => r := "01001011011100001010111110011110111";
      when 3450 => r := "01001011011000001010111101010011100";
      when 3451 => r := "01001011011000001010111100001000000";
      when 3452 => r := "01001011010100001010111010111100100";
      when 3453 => r := "01001011010100001010111001110001010";
      when 3454 => r := "01001011010100001010111000100110000";
      when 3455 => r := "01001011010100001010110111011010101";
      when 3456 => r := "01001011010000001010110110001111001";
      when 3457 => r := "01001011010000001010110101000011111";
      when 3458 => r := "01001011001100001010110011111000101";
      when 3459 => r := "01001011001100001010110010101101100";
      when 3460 => r := "01001011001100001010110001100010000";
      when 3461 => r := "01001011001100001010110000010110111";
      when 3462 => r := "01001011001000001010101111001011101";
      when 3463 => r := "01001011001000001010101110000000100";
      when 3464 => r := "01001011001000001010101100110101100";
      when 3465 => r := "01001011001000001010101011101010011";
      when 3466 => r := "01001011000100001010101010011111010";
      when 3467 => r := "01001011000100001010101001010100001";
      when 3468 => r := "01001011000000001010101000001001000";
      when 3469 => r := "01001011000000001010100110111110000";
      when 3470 => r := "01001011000000001010100101110010110";
      when 3471 => r := "01001011000000001010100100100111110";
      when 3472 => r := "01001010111100001010100011011100110";
      when 3473 => r := "01001010111100001010100010010001110";
      when 3474 => r := "01001010111000001010100001000110111";
      when 3475 => r := "01001010111000001010011111111100000";
      when 3476 => r := "01001010111000001010011110110001000";
      when 3477 => r := "01001010111000001010011101100110001";
      when 3478 => r := "01001010110100001010011100011011010";
      when 3479 => r := "01001010110100001010011011010000011";
      when 3480 => r := "01001010110000001010011010000101101";
      when 3481 => r := "01001010110000001010011000111010110";
      when 3482 => r := "01001010110000001010010111101111111";
      when 3483 => r := "01001010110000001010010110100101001";
      when 3484 => r := "01001010101100001010010101011010011";
      when 3485 => r := "01001010101100001010010100001111101";
      when 3486 => r := "01001010101100001010010011000101000";
      when 3487 => r := "01001010101100001010010001111010010";
      when 3488 => r := "01001010101000001010010000101111101";
      when 3489 => r := "01001010101000001010001111100101000";
      when 3490 => r := "01001010100100001010001110011010010";
      when 3491 => r := "01001010100100001010001101001111110";
      when 3492 => r := "01001010100100001010001100000101001";
      when 3493 => r := "01001010100100001010001010111010100";
      when 3494 => r := "01001010100000001010001001101111111";
      when 3495 => r := "01001010100000001010001000100101011";
      when 3496 => r := "01001010011100001010000111011010111";
      when 3497 => r := "01001010011100001010000110010000011";
      when 3498 => r := "01001010011100001010000101000101111";
      when 3499 => r := "01001010011100001010000011111011011";
      when 3500 => r := "01001010011000001010000010110000111";
      when 3501 => r := "01001010011000001010000001100110100";
      when 3502 => r := "01001010011000001010000000011100001";
      when 3503 => r := "01001010011000001001111111010001110";
      when 3504 => r := "01001010010100001001111110000111011";
      when 3505 => r := "01001010010100001001111100111101000";
      when 3506 => r := "01001010010000001001111011110010100";
      when 3507 => r := "01001010010000001001111010101000010";
      when 3508 => r := "01001010010000001001111001011110001";
      when 3509 => r := "01001010010000001001111000010011110";
      when 3510 => r := "01001010001100001001110111001001100";
      when 3511 => r := "01001010001100001001110101111111010";
      when 3512 => r := "01001010001000001001110100110101000";
      when 3513 => r := "01001010001000001001110011101010111";
      when 3514 => r := "01001010001000001001110010100000110";
      when 3515 => r := "01001010001000001001110001010110101";
      when 3516 => r := "01001010000100001001110000001100011";
      when 3517 => r := "01001010000100001001101111000010010";
      when 3518 => r := "01001010000100001001101101111000010";
      when 3519 => r := "01001010000100001001101100101110001";
      when 3520 => r := "01001010000000001001101011100100001";
      when 3521 => r := "01001010000000001001101010011010000";
      when 3522 => r := "01001001111100001001101001001111111";
      when 3523 => r := "01001001111100001001101000000101111";
      when 3524 => r := "01001001111100001001100110111011111";
      when 3525 => r := "01001001111100001001100101110010000";
      when 3526 => r := "01001001111000001001100100101000010";
      when 3527 => r := "01001001111000001001100011011110011";
      when 3528 => r := "01001001110100001001100010010100011";
      when 3529 => r := "01001001110100001001100001001010100";
      when 3530 => r := "01001001110100001001100000000000100";
      when 3531 => r := "01001001110100001001011110110110110";
      when 3532 => r := "01001001110000001001011101101101000";
      when 3533 => r := "01001001110000001001011100100011010";
      when 3534 => r := "01001001110000001001011011011001011";
      when 3535 => r := "01001001110000001001011010001111101";
      when 3536 => r := "01001001101100001001011001000101111";
      when 3537 => r := "01001001101100001001010111111100001";
      when 3538 => r := "01001001101000001001010110110010010";
      when 3539 => r := "01001001101000001001010101101000101";
      when 3540 => r := "01001001101000001001010100011111000";
      when 3541 => r := "01001001101000001001010011010101011";
      when 3542 => r := "01001001100100001001010010001011110";
      when 3543 => r := "01001001100100001001010001000010001";
      when 3544 => r := "01001001100100001001001111111000100";
      when 3545 => r := "01001001100100001001001110101111000";
      when 3546 => r := "01001001100000001001001101100101011";
      when 3547 => r := "01001001100000001001001100011011111";
      when 3548 => r := "01001001011100001001001011010010100";
      when 3549 => r := "01001001011100001001001010001001000";
      when 3550 => r := "01001001011100001001001000111111011";
      when 3551 => r := "01001001011100001001000111110110000";
      when 3552 => r := "01001001011000001001000110101100011";
      when 3553 => r := "01001001011000001001000101100011000";
      when 3554 => r := "01001001010100001001000100011001110";
      when 3555 => r := "01001001010100001001000011010000011";
      when 3556 => r := "01001001010100001001000010000111001";
      when 3557 => r := "01001001010100001001000000111101110";
      when 3558 => r := "01001001010000001000111111110100010";
      when 3559 => r := "01001001010000001000111110101011000";
      when 3560 => r := "01001001010000001000111101100001101";
      when 3561 => r := "01001001010000001000111100011000011";
      when 3562 => r := "01001001001100001000111011001111010";
      when 3563 => r := "01001001001100001000111010000110000";
      when 3564 => r := "01001001001000001000111000111100101";
      when 3565 => r := "01001001001000001000110111110011100";
      when 3566 => r := "01001001001000001000110110101010010";
      when 3567 => r := "01001001001000001000110101100001001";
      when 3568 => r := "01001001000100001000110100011000001";
      when 3569 => r := "01001001000100001000110011001111000";
      when 3570 => r := "01001001000100001000110010000101110";
      when 3571 => r := "01001001000100001000110000111100110";
      when 3572 => r := "01001001000000001000101111110011110";
      when 3573 => r := "01001001000000001000101110101010110";
      when 3574 => r := "01001000111100001000101101100001110";
      when 3575 => r := "01001000111100001000101100011000110";
      when 3576 => r := "01001000111100001000101011001111110";
      when 3577 => r := "01001000111100001000101010000110111";
      when 3578 => r := "01001000111000001000101000111101110";
      when 3579 => r := "01001000111000001000100111110100111";
      when 3580 => r := "01001000110100001000100110101100000";
      when 3581 => r := "01001000110100001000100101100011001";
      when 3582 => r := "01001000110100001000100100011010010";
      when 3583 => r := "01001000110100001000100011010001011";
      when 3584 => r := "01001000110000001000100010001000101";
      when 3585 => r := "01001000110000001000100000111111110";
      when 3586 => r := "01001000110000001000011111110111000";
      when 3587 => r := "01001000110000001000011110101110010";
      when 3588 => r := "01001000101100001000011101100101100";
      when 3589 => r := "01001000101100001000011100011100110";
      when 3590 => r := "01001000101000001000011011010100000";
      when 3591 => r := "01001000101000001000011010001011010";
      when 3592 => r := "01001000101000001000011001000010100";
      when 3593 => r := "01001000101000001000010111111001111";
      when 3594 => r := "01001000100100001000010110110001011";
      when 3595 => r := "01001000100100001000010101101000110";
      when 3596 => r := "01001000100100001000010100100000010";
      when 3597 => r := "01001000100100001000010011010111101";
      when 3598 => r := "01001000100000001000010010001111000";
      when 3599 => r := "01001000100000001000010001000110100";
      when 3600 => r := "01001000011100001000001111111101111";
      when 3601 => r := "01001000011100001000001110110101011";
      when 3602 => r := "01001000011100001000001101101100110";
      when 3603 => r := "01001000011100001000001100100100011";
      when 3604 => r := "01001000011000001000001011011100000";
      when 3605 => r := "01001000011000001000001010010011100";
      when 3606 => r := "01001000011000001000001001001011001";
      when 3607 => r := "01001000011000001000001000000010110";
      when 3608 => r := "01001000010100001000000110111010011";
      when 3609 => r := "01001000010100001000000101110010000";
      when 3610 => r := "01001000010000001000000100101001110";
      when 3611 => r := "01001000010000001000000011100001100";
      when 3612 => r := "01001000010000001000000010011001000";
      when 3613 => r := "01001000010000001000000001010000110";
      when 3614 => r := "01001000001100001000000000001000100";
      when 3615 => r := "01001000001100000111111111000000010";
      when 3616 => r := "01001000001100000111111101111000000";
      when 3617 => r := "01001000001100000111111100101111110";
      when 3618 => r := "01001000001000000111111011100111110";
      when 3619 => r := "01001000001000000111111010011111100";
      when 3620 => r := "01001000000100000111111001010111011";
      when 3621 => r := "01001000000100000111111000001111010";
      when 3622 => r := "01001000000100000111110111000111001";
      when 3623 => r := "01001000000100000111110101111111001";
      when 3624 => r := "01001000000000000111110100110111000";
      when 3625 => r := "01001000000000000111110011101110111";
      when 3626 => r := "01001000000000000111110010100110110";
      when 3627 => r := "01001000000000000111110001011110110";
      when 3628 => r := "01000111111100000111110000010110111";
      when 3629 => r := "01000111111100000111101111001111000";
      when 3630 => r := "01000111111000000111101110000111000";
      when 3631 => r := "01000111111000000111101100111111000";
      when 3632 => r := "01000111111000000111101011110111000";
      when 3633 => r := "01000111111000000111101010101111001";
      when 3634 => r := "01000111110100000111101001100111010";
      when 3635 => r := "01000111110100000111101000011111011";
      when 3636 => r := "01000111110100000111100111010111101";
      when 3637 => r := "01000111110100000111100110001111110";
      when 3638 => r := "01000111110000000111100101000111110";
      when 3639 => r := "01000111110000000111100100000000000";
      when 3640 => r := "01000111101100000111100010111000010";
      when 3641 => r := "01000111101100000111100001110000101";
      when 3642 => r := "01000111101100000111100000101000111";
      when 3643 => r := "01000111101100000111011111100001001";
      when 3644 => r := "01000111101000000111011110011001011";
      when 3645 => r := "01000111101000000111011101010001110";
      when 3646 => r := "01000111101000000111011100001010001";
      when 3647 => r := "01000111101000000111011011000010100";
      when 3648 => r := "01000111100100000111011001111010110";
      when 3649 => r := "01000111100100000111011000110011001";
      when 3650 => r := "01000111100100000111010111101011100";
      when 3651 => r := "01000111100100000111010110100100000";
      when 3652 => r := "01000111100000000111010101011100100";
      when 3653 => r := "01000111100000000111010100010101000";
      when 3654 => r := "01000111011100000111010011001101011";
      when 3655 => r := "01000111011100000111010010000110000";
      when 3656 => r := "01000111011100000111010000111110100";
      when 3657 => r := "01000111011100000111001111110111000";
      when 3658 => r := "01000111011000000111001110101111011";
      when 3659 => r := "01000111011000000111001101101000000";
      when 3660 => r := "01000111011000000111001100100000101";
      when 3661 => r := "01000111011000000111001011011001010";
      when 3662 => r := "01000111010100000111001010010010000";
      when 3663 => r := "01000111010100000111001001001010101";
      when 3664 => r := "01000111010000000111001000000011010";
      when 3665 => r := "01000111010000000111000110111100000";
      when 3666 => r := "01000111010000000111000101110100101";
      when 3667 => r := "01000111010000000111000100101101011";
      when 3668 => r := "01000111001100000111000011100110000";
      when 3669 => r := "01000111001100000111000010011110110";
      when 3670 => r := "01000111001100000111000001010111100";
      when 3671 => r := "01000111001100000111000000010000010";
      when 3672 => r := "01000111001000000110111111001001001";
      when 3673 => r := "01000111001000000110111110000010000";
      when 3674 => r := "01000111000100000110111100111010110";
      when 3675 => r := "01000111000100000110111011110011101";
      when 3676 => r := "01000111000100000110111010101100101";
      when 3677 => r := "01000111000100000110111001100101100";
      when 3678 => r := "01000111000000000110111000011110101";
      when 3679 => r := "01000111000000000110110111010111100";
      when 3680 => r := "01000111000000000110110110010000011";
      when 3681 => r := "01000111000000000110110101001001011";
      when 3682 => r := "01000110111100000110110100000010010";
      when 3683 => r := "01000110111100000110110010111011010";
      when 3684 => r := "01000110111100000110110001110100011";
      when 3685 => r := "01000110111100000110110000101101100";
      when 3686 => r := "01000110111000000110101111100110101";
      when 3687 => r := "01000110111000000110101110011111110";
      when 3688 => r := "01000110110100000110101101011000110";
      when 3689 => r := "01000110110100000110101100010001111";
      when 3690 => r := "01000110110100000110101011001010111";
      when 3691 => r := "01000110110100000110101010000100001";
      when 3692 => r := "01000110110000000110101000111101011";
      when 3693 => r := "01000110110000000110100111110110101";
      when 3694 => r := "01000110110000000110100110101111101";
      when 3695 => r := "01000110110000000110100101101000111";
      when 3696 => r := "01000110101100000110100100100010010";
      when 3697 => r := "01000110101100000110100011011011100";
      when 3698 => r := "01000110101000000110100010010100110";
      when 3699 => r := "01000110101000000110100001001110001";
      when 3700 => r := "01000110101000000110100000000111011";
      when 3701 => r := "01000110101000000110011111000000110";
      when 3702 => r := "01000110100100000110011101111010010";
      when 3703 => r := "01000110100100000110011100110011101";
      when 3704 => r := "01000110100100000110011011101100111";
      when 3705 => r := "01000110100100000110011010100110010";
      when 3706 => r := "01000110100000000110011001011111110";
      when 3707 => r := "01000110100000000110011000011001001";
      when 3708 => r := "01000110100000000110010111010010100";
      when 3709 => r := "01000110100000000110010110001100000";
      when 3710 => r := "01000110011100000110010101000101100";
      when 3711 => r := "01000110011100000110010011111111001";
      when 3712 => r := "01000110011000000110010010111000101";
      when 3713 => r := "01000110011000000110010001110010010";
      when 3714 => r := "01000110011000000110010000101011110";
      when 3715 => r := "01000110011000000110001111100101011";
      when 3716 => r := "01000110010100000110001110011111000";
      when 3717 => r := "01000110010100000110001101011000101";
      when 3718 => r := "01000110010100000110001100010010010";
      when 3719 => r := "01000110010100000110001011001100000";
      when 3720 => r := "01000110010000000110001010000101110";
      when 3721 => r := "01000110010000000110001000111111100";
      when 3722 => r := "01000110010000000110000111111001001";
      when 3723 => r := "01000110010000000110000110110010111";
      when 3724 => r := "01000110001100000110000101101100100";
      when 3725 => r := "01000110001100000110000100100110011";
      when 3726 => r := "01000110001000000110000011100000001";
      when 3727 => r := "01000110001000000110000010011010000";
      when 3728 => r := "01000110001000000110000001010011101";
      when 3729 => r := "01000110001000000110000000001101100";
      when 3730 => r := "01000110000100000101111111000111011";
      when 3731 => r := "01000110000100000101111110000001010";
      when 3732 => r := "01000110000100000101111100111011010";
      when 3733 => r := "01000110000100000101111011110101010";
      when 3734 => r := "01000110000000000101111010101111001";
      when 3735 => r := "01000110000000000101111001101001001";
      when 3736 => r := "01000110000000000101111000100011000";
      when 3737 => r := "01000110000000000101110111011101000";
      when 3738 => r := "01000101111100000101110110010111001";
      when 3739 => r := "01000101111100000101110101010001010";
      when 3740 => r := "01000101111000000101110100001011001";
      when 3741 => r := "01000101111000000101110011000101010";
      when 3742 => r := "01000101111000000101110001111111001";
      when 3743 => r := "01000101111000000101110000111001010";
      when 3744 => r := "01000101110100000101101111110011100";
      when 3745 => r := "01000101110100000101101110101101101";
      when 3746 => r := "01000101110100000101101101100111101";
      when 3747 => r := "01000101110100000101101100100001111";
      when 3748 => r := "01000101110000000101101011011100001";
      when 3749 => r := "01000101110000000101101010010110011";
      when 3750 => r := "01000101110000000101101001010000101";
      when 3751 => r := "01000101110000000101101000001010111";
      when 3752 => r := "01000101101100000101100111000101000";
      when 3753 => r := "01000101101100000101100101111111010";
      when 3754 => r := "01000101101000000101100100111001110";
      when 3755 => r := "01000101101000000101100011110100000";
      when 3756 => r := "01000101101000000101100010101110010";
      when 3757 => r := "01000101101000000101100001101000101";
      when 3758 => r := "01000101100100000101100000100011000";
      when 3759 => r := "01000101100100000101011111011101100";
      when 3760 => r := "01000101100100000101011110010111110";
      when 3761 => r := "01000101100100000101011101010010010";
      when 3762 => r := "01000101100000000101011100001100100";
      when 3763 => r := "01000101100000000101011011000111000";
      when 3764 => r := "01000101100000000101011010000001100";
      when 3765 => r := "01000101100000000101011000111011111";
      when 3766 => r := "01000101011100000101010111110110100";
      when 3767 => r := "01000101011100000101010110110001000";
      when 3768 => r := "01000101011000000101010101101011100";
      when 3769 => r := "01000101011000000101010100100110001";
      when 3770 => r := "01000101011000000101010011100000101";
      when 3771 => r := "01000101011000000101010010011011010";
      when 3772 => r := "01000101010100000101010001010110000";
      when 3773 => r := "01000101010100000101010000010000101";
      when 3774 => r := "01000101010100000101001111001011010";
      when 3775 => r := "01000101010100000101001110000110000";
      when 3776 => r := "01000101010000000101001101000000100";
      when 3777 => r := "01000101010000000101001011111011001";
      when 3778 => r := "01000101010000000101001010110110000";
      when 3779 => r := "01000101010000000101001001110000110";
      when 3780 => r := "01000101001100000101001000101011101";
      when 3781 => r := "01000101001100000101000111100110011";
      when 3782 => r := "01000101001000000101000110100001000";
      when 3783 => r := "01000101001000000101000101011011111";
      when 3784 => r := "01000101001000000101000100010110101";
      when 3785 => r := "01000101001000000101000011010001100";
      when 3786 => r := "01000101000100000101000010001100010";
      when 3787 => r := "01000101000100000101000001000111001";
      when 3788 => r := "01000101000100000101000000000010001";
      when 3789 => r := "01000101000100000100111110111101000";
      when 3790 => r := "01000101000000000100111101110111110";
      when 3791 => r := "01000101000000000100111100110010110";
      when 3792 => r := "01000101000000000100111011101101111";
      when 3793 => r := "01000101000000000100111010101000111";
      when 3794 => r := "01000100111100000100111001100011111";
      when 3795 => r := "01000100111100000100111000011111000";
      when 3796 => r := "01000100111100000100110111011001110";
      when 3797 => r := "01000100111100000100110110010100111";
      when 3798 => r := "01000100111000000100110101010000000";
      when 3799 => r := "01000100111000000100110100001011001";
      when 3800 => r := "01000100110100000100110011000110010";
      when 3801 => r := "01000100110100000100110010000001011";
      when 3802 => r := "01000100110100000100110000111100100";
      when 3803 => r := "01000100110100000100101111110111101";
      when 3804 => r := "01000100110000000100101110110010110";
      when 3805 => r := "01000100110000000100101101101110000";
      when 3806 => r := "01000100110000000100101100101001001";
      when 3807 => r := "01000100110000000100101011100100011";
      when 3808 => r := "01000100101100000100101010011111101";
      when 3809 => r := "01000100101100000100101001011010111";
      when 3810 => r := "01000100101100000100101000010110001";
      when 3811 => r := "01000100101100000100100111010001011";
      when 3812 => r := "01000100101000000100100110001100110";
      when 3813 => r := "01000100101000000100100101001000001";
      when 3814 => r := "01000100101000000100100100000011100";
      when 3815 => r := "01000100101000000100100010111110111";
      when 3816 => r := "01000100100100000100100001111010001";
      when 3817 => r := "01000100100100000100100000110101101";
      when 3818 => r := "01000100100000000100011111110001000";
      when 3819 => r := "01000100100000000100011110101100100";
      when 3820 => r := "01000100100000000100011101100111111";
      when 3821 => r := "01000100100000000100011100100011011";
      when 3822 => r := "01000100011100000100011011011110111";
      when 3823 => r := "01000100011100000100011010011010011";
      when 3824 => r := "01000100011100000100011001010101111";
      when 3825 => r := "01000100011100000100011000010001011";
      when 3826 => r := "01000100011000000100010111001101000";
      when 3827 => r := "01000100011000000100010110001000100";
      when 3828 => r := "01000100011000000100010101000100001";
      when 3829 => r := "01000100011000000100010011111111110";
      when 3830 => r := "01000100010100000100010010111011010";
      when 3831 => r := "01000100010100000100010001110110111";
      when 3832 => r := "01000100010100000100010000110010101";
      when 3833 => r := "01000100010100000100001111101110011";
      when 3834 => r := "01000100010000000100001110101010001";
      when 3835 => r := "01000100010000000100001101100101110";
      when 3836 => r := "01000100001100000100001100100001100";
      when 3837 => r := "01000100001100000100001011011101010";
      when 3838 => r := "01000100001100000100001010011000111";
      when 3839 => r := "01000100001100000100001001010100101";
      when 3840 => r := "01000100001000000100001000010000101";
      when 3841 => r := "01000100001000000100000111001100100";
      when 3842 => r := "01000100001000000100000110001000001";
      when 3843 => r := "01000100001000000100000101000100000";
      when 3844 => r := "01000100000100000100000100000000000";
      when 3845 => r := "01000100000100000100000010111011111";
      when 3846 => r := "01000100000100000100000001110111110";
      when 3847 => r := "01000100000100000100000000110011110";
      when 3848 => r := "01000100000000000011111111101111100";
      when 3849 => r := "01000100000000000011111110101011100";
      when 3850 => r := "01000100000000000011111101100111011";
      when 3851 => r := "01000100000000000011111100100011011";
      when 3852 => r := "01000011111100000011111011011111100";
      when 3853 => r := "01000011111100000011111010011011100";
      when 3854 => r := "01000011111100000011111001010111100";
      when 3855 => r := "01000011111100000011111000010011100";
      when 3856 => r := "01000011111000000011110111001111101";
      when 3857 => r := "01000011111000000011110110001011110";
      when 3858 => r := "01000011110100000011110101000111110";
      when 3859 => r := "01000011110100000011110100000011111";
      when 3860 => r := "01000011110100000011110011000000000";
      when 3861 => r := "01000011110100000011110001111100010";
      when 3862 => r := "01000011110000000011110000111000011";
      when 3863 => r := "01000011110000000011101111110100101";
      when 3864 => r := "01000011110000000011101110110000111";
      when 3865 => r := "01000011110000000011101101101101001";
      when 3866 => r := "01000011101100000011101100101001001";
      when 3867 => r := "01000011101100000011101011100101011";
      when 3868 => r := "01000011101100000011101010100001110";
      when 3869 => r := "01000011101100000011101001011110001";
      when 3870 => r := "01000011101000000011101000011010010";
      when 3871 => r := "01000011101000000011100111010110101";
      when 3872 => r := "01000011101000000011100110010011001";
      when 3873 => r := "01000011101000000011100101001111100";
      when 3874 => r := "01000011100100000011100100001011111";
      when 3875 => r := "01000011100100000011100011001000010";
      when 3876 => r := "01000011100100000011100010000100101";
      when 3877 => r := "01000011100100000011100001000001000";
      when 3878 => r := "01000011100000000011011111111101011";
      when 3879 => r := "01000011100000000011011110111001111";
      when 3880 => r := "01000011011100000011011101110110011";
      when 3881 => r := "01000011011100000011011100110010111";
      when 3882 => r := "01000011011100000011011011101111100";
      when 3883 => r := "01000011011100000011011010101100000";
      when 3884 => r := "01000011011000000011011001101000100";
      when 3885 => r := "01000011011000000011011000100101001";
      when 3886 => r := "01000011011000000011010111100001101";
      when 3887 => r := "01000011011000000011010110011110010";
      when 3888 => r := "01000011010100000011010101011010110";
      when 3889 => r := "01000011010100000011010100010111100";
      when 3890 => r := "01000011010100000011010011010100000";
      when 3891 => r := "01000011010100000011010010010000101";
      when 3892 => r := "01000011010000000011010001001101011";
      when 3893 => r := "01000011010000000011010000001010000";
      when 3894 => r := "01000011010000000011001111000110111";
      when 3895 => r := "01000011010000000011001110000011101";
      when 3896 => r := "01000011001100000011001101000000010";
      when 3897 => r := "01000011001100000011001011111101000";
      when 3898 => r := "01000011001100000011001010111001111";
      when 3899 => r := "01000011001100000011001001110110110";
      when 3900 => r := "01000011001000000011001000110011100";
      when 3901 => r := "01000011001000000011000111110000011";
      when 3902 => r := "01000011001000000011000110101101010";
      when 3903 => r := "01000011001000000011000101101010001";
      when 3904 => r := "01000011000100000011000100100110111";
      when 3905 => r := "01000011000100000011000011100011111";
      when 3906 => r := "01000011000000000011000010100000101";
      when 3907 => r := "01000011000000000011000001011101101";
      when 3908 => r := "01000011000000000011000000011010110";
      when 3909 => r := "01000011000000000010111111010111110";
      when 3910 => r := "01000010111100000010111110010100101";
      when 3911 => r := "01000010111100000010111101010001101";
      when 3912 => r := "01000010111100000010111100001110101";
      when 3913 => r := "01000010111100000010111011001011110";
      when 3914 => r := "01000010111000000010111010001000110";
      when 3915 => r := "01000010111000000010111001000101110";
      when 3916 => r := "01000010111000000010111000000010111";
      when 3917 => r := "01000010111000000010110111000000000";
      when 3918 => r := "01000010110100000010110101111101001";
      when 3919 => r := "01000010110100000010110100111010010";
      when 3920 => r := "01000010110100000010110011110111011";
      when 3921 => r := "01000010110100000010110010110100100";
      when 3922 => r := "01000010110000000010110001110001110";
      when 3923 => r := "01000010110000000010110000101110111";
      when 3924 => r := "01000010110000000010101111101100001";
      when 3925 => r := "01000010110000000010101110101001011";
      when 3926 => r := "01000010101100000010101101100110101";
      when 3927 => r := "01000010101100000010101100100011111";
      when 3928 => r := "01000010101100000010101011100001001";
      when 3929 => r := "01000010101100000010101010011110100";
      when 3930 => r := "01000010101000000010101001011011111";
      when 3931 => r := "01000010101000000010101000011001010";
      when 3932 => r := "01000010100100000010100111010110100";
      when 3933 => r := "01000010100100000010100110010011111";
      when 3934 => r := "01000010100100000010100101010001010";
      when 3935 => r := "01000010100100000010100100001110110";
      when 3936 => r := "01000010100000000010100011001100000";
      when 3937 => r := "01000010100000000010100010001001100";
      when 3938 => r := "01000010100000000010100001000110110";
      when 3939 => r := "01000010100000000010100000000100010";
      when 3940 => r := "01000010011100000010011111000001111";
      when 3941 => r := "01000010011100000010011101111111011";
      when 3942 => r := "01000010011100000010011100111100110";
      when 3943 => r := "01000010011100000010011011111010011";
      when 3944 => r := "01000010011000000010011010111000000";
      when 3945 => r := "01000010011000000010011001110101100";
      when 3946 => r := "01000010011000000010011000110011000";
      when 3947 => r := "01000010011000000010010111110000101";
      when 3948 => r := "01000010010100000010010110101110011";
      when 3949 => r := "01000010010100000010010101101100000";
      when 3950 => r := "01000010010100000010010100101001100";
      when 3951 => r := "01000010010100000010010011100111001";
      when 3952 => r := "01000010010000000010010010100101000";
      when 3953 => r := "01000010010000000010010001100010101";
      when 3954 => r := "01000010010000000010010000100000010";
      when 3955 => r := "01000010010000000010001111011110000";
      when 3956 => r := "01000010001100000010001110011011111";
      when 3957 => r := "01000010001100000010001101011001101";
      when 3958 => r := "01000010001100000010001100010111100";
      when 3959 => r := "01000010001100000010001011010101010";
      when 3960 => r := "01000010001000000010001010010011000";
      when 3961 => r := "01000010001000000010001001010000111";
      when 3962 => r := "01000010001000000010001000001110100";
      when 3963 => r := "01000010001000000010000111001100011";
      when 3964 => r := "01000010000100000010000110001010011";
      when 3965 => r := "01000010000100000010000101001000010";
      when 3966 => r := "01000010000100000010000100000110001";
      when 3967 => r := "01000010000100000010000011000100001";
      when 3968 => r := "01000010000000000010000010000010000";
      when 3969 => r := "01000010000000000010000001000000000";
      when 3970 => r := "01000001111100000001111111111101111";
      when 3971 => r := "01000001111100000001111110111100000";
      when 3972 => r := "01000001111100000001111101111001111";
      when 3973 => r := "01000001111100000001111100110111111";
      when 3974 => r := "01000001111000000001111011110110000";
      when 3975 => r := "01000001111000000001111010110100000";
      when 3976 => r := "01000001111000000001111001110010010";
      when 3977 => r := "01000001111000000001111000110000011";
      when 3978 => r := "01000001110100000001110111101110011";
      when 3979 => r := "01000001110100000001110110101100100";
      when 3980 => r := "01000001110100000001110101101010101";
      when 3981 => r := "01000001110100000001110100101000110";
      when 3982 => r := "01000001110000000001110011100110111";
      when 3983 => r := "01000001110000000001110010100101001";
      when 3984 => r := "01000001110000000001110001100011011";
      when 3985 => r := "01000001110000000001110000100001101";
      when 3986 => r := "01000001101100000001101111011111110";
      when 3987 => r := "01000001101100000001101110011110001";
      when 3988 => r := "01000001101100000001101101011100011";
      when 3989 => r := "01000001101100000001101100011010101";
      when 3990 => r := "01000001101000000001101011011001000";
      when 3991 => r := "01000001101000000001101010010111010";
      when 3992 => r := "01000001101000000001101001010101101";
      when 3993 => r := "01000001101000000001101000010100000";
      when 3994 => r := "01000001100100000001100111010010011";
      when 3995 => r := "01000001100100000001100110010000110";
      when 3996 => r := "01000001100100000001100101001111001";
      when 3997 => r := "01000001100100000001100100001101100";
      when 3998 => r := "01000001100000000001100011001100000";
      when 3999 => r := "01000001100000000001100010001010100";
      when 4000 => r := "01000001100000000001100001001000111";
      when 4001 => r := "01000001100000000001100000000111011";
      when 4002 => r := "01000001011100000001011111000101110";
      when 4003 => r := "01000001011100000001011110000100011";
      when 4004 => r := "01000001011100000001011101000010110";
      when 4005 => r := "01000001011100000001011100000001011";
      when 4006 => r := "01000001011000000001011011000000000";
      when 4007 => r := "01000001011000000001011001111110101";
      when 4008 => r := "01000001011000000001011000111101001";
      when 4009 => r := "01000001011000000001010111111011110";
      when 4010 => r := "01000001010100000001010110111010100";
      when 4011 => r := "01000001010100000001010101111001001";
      when 4012 => r := "01000001010100000001010100110111110";
      when 4013 => r := "01000001010100000001010011110110011";
      when 4014 => r := "01000001010000000001010010110101000";
      when 4015 => r := "01000001010000000001010001110011110";
      when 4016 => r := "01000001010000000001010000110010011";
      when 4017 => r := "01000001010000000001001111110001001";
      when 4018 => r := "01000001001100000001001110110000000";
      when 4019 => r := "01000001001100000001001101101110110";
      when 4020 => r := "01000001001100000001001100101101101";
      when 4021 => r := "01000001001100000001001011101100011";
      when 4022 => r := "01000001001000000001001010101011001";
      when 4023 => r := "01000001001000000001001001101010000";
      when 4024 => r := "01000001000100000001001000101000110";
      when 4025 => r := "01000001000100000001000111100111101";
      when 4026 => r := "01000001000100000001000110100110101";
      when 4027 => r := "01000001000100000001000101100101100";
      when 4028 => r := "01000001000000000001000100100100100";
      when 4029 => r := "01000001000000000001000011100011011";
      when 4030 => r := "01000001000000000001000010100010010";
      when 4031 => r := "01000001000000000001000001100001010";
      when 4032 => r := "01000000111100000001000000100000010";
      when 4033 => r := "01000000111100000000111111011111010";
      when 4034 => r := "01000000111100000000111110011110010";
      when 4035 => r := "01000000111100000000111101011101010";
      when 4036 => r := "01000000111000000000111100011100011";
      when 4037 => r := "01000000111000000000111011011011011";
      when 4038 => r := "01000000111000000000111010011010100";
      when 4039 => r := "01000000111000000000111001011001101";
      when 4040 => r := "01000000110100000000111000011000110";
      when 4041 => r := "01000000110100000000110111010111111";
      when 4042 => r := "01000000110100000000110110010111000";
      when 4043 => r := "01000000110100000000110101010110001";
      when 4044 => r := "01000000110000000000110100010101011";
      when 4045 => r := "01000000110000000000110011010100101";
      when 4046 => r := "01000000110000000000110010010011101";
      when 4047 => r := "01000000110000000000110001010010111";
      when 4048 => r := "01000000101100000000110000010010001";
      when 4049 => r := "01000000101100000000101111010001011";
      when 4050 => r := "01000000101100000000101110010000110";
      when 4051 => r := "01000000101100000000101101010000000";
      when 4052 => r := "01000000101000000000101100001111011";
      when 4053 => r := "01000000101000000000101011001110101";
      when 4054 => r := "01000000101000000000101010001101111";
      when 4055 => r := "01000000101000000000101001001101010";
      when 4056 => r := "01000000100100000000101000001100110";
      when 4057 => r := "01000000100100000000100111001100001";
      when 4058 => r := "01000000100100000000100110001011011";
      when 4059 => r := "01000000100100000000100101001010110";
      when 4060 => r := "01000000100000000000100100001010001";
      when 4061 => r := "01000000100000000000100011001001100";
      when 4062 => r := "01000000100000000000100010001001000";
      when 4063 => r := "01000000100000000000100001001000100";
      when 4064 => r := "01000000011100000000100000001000001";
      when 4065 => r := "01000000011100000000011111000111101";
      when 4066 => r := "01000000011100000000011110000111000";
      when 4067 => r := "01000000011100000000011101000110101";
      when 4068 => r := "01000000011000000000011100000110010";
      when 4069 => r := "01000000011000000000011011000101110";
      when 4070 => r := "01000000011000000000011010000101011";
      when 4071 => r := "01000000011000000000011001000101000";
      when 4072 => r := "01000000010100000000011000000100100";
      when 4073 => r := "01000000010100000000010111000100001";
      when 4074 => r := "01000000010100000000010110000011110";
      when 4075 => r := "01000000010100000000010101000011100";
      when 4076 => r := "01000000010000000000010100000011010";
      when 4077 => r := "01000000010000000000010011000011000";
      when 4078 => r := "01000000010000000000010010000010101";
      when 4079 => r := "01000000010000000000010001000010011";
      when 4080 => r := "01000000001100000000010000000010000";
      when 4081 => r := "01000000001100000000001111000001110";
      when 4082 => r := "01000000001100000000001110000001100";
      when 4083 => r := "01000000001100000000001101000001011";
      when 4084 => r := "01000000001000000000001100000001001";
      when 4085 => r := "01000000001000000000001011000001000";
      when 4086 => r := "01000000001000000000001010000000110";
      when 4087 => r := "01000000001000000000001001000000101";
      when 4088 => r := "01000000000100000000001000000000100";
      when 4089 => r := "01000000000100000000000111000000011";
      when 4090 => r := "01000000000100000000000110000000010";
      when 4091 => r := "01000000000100000000000101000000010";
      when 4092 => r := "01000000000000000000000100000000001";
      when 4093 => r := "01000000000000000000000011000000001";
      when 4094 => r := "01000000000000000000000010000000000";
      when 4095 => r := "01000000000000000000000001000000000";
      when others => r := (others => '0');
    end case;
    return r;
  end table;

  signal ret : std_logic_vector (31 downto 0) := (others => '0');
  signal sign : std_logic := '0';
  signal expr : std_logic_vector (7 downto 0) := (others => '0');
  signal expr2 : std_logic_vector (7 downto 0) := (others => '0');
  signal key : std_logic_vector (11 downto 0) := (others => '0');
  signal i_mantissa : std_logic_vector (22 downto 0) := (others => '0');
  signal o_mantissa : std_logic_vector (22 downto 0) := (others => '0');
  signal l_b : std_logic_vector (10 downto 0) := (others => '0');
  signal HL : std_logic_vector (22 downto 0) := (others => '0');
  signal raw_ret : std_logic_vector (34 downto 0) := (others => '0');
  signal ret_a : std_logic_vector (11 downto 0) := (others => '0');
  signal ret_b : std_logic_vector (22 downto 0) := (others => '0');
  signal mul : std_logic_vector (10 downto 0) := (others => '0');
begin -- architecture rtl

  with i_mantissa select
    ret <=
    sign & expr2 & "00000000000000000000000" when "00000000000000000000000",
    sign & expr & o_mantissa (21 downto 0) & '0' when others;

  sign <= a (31);
  expr <= 126 + 127 - a (30 downto 23);
  expr2 <= 127 + 127 - a (30 downto 23);
  i_mantissa <= a (22 downto 0);
  l_b <= a (10 downto 0);
  key <= a (22 downto 11);
  raw_ret <= table (key);
  ret_a <= raw_ret (34 downto 23);
  ret_b <= raw_ret (22 downto 0);
  HL <= ret_a * l_b;
  mul <= HL (22 downto 12);
  o_mantissa <= "00000000000000000000000" + ((ret_b - mul));

  -- purpose: set ret -> Q
  -- type : combinational
  -- inputs : CLK
  -- outputs: Q
  set_loop: process (CLK) is
  begin -- process set_loop
    if rising_edge (CLK) then
      Q <= ret;
    end if;
  end process set_loop;

end architecture rtl;
