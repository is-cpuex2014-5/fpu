library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity fsqrt is  
  port (
    A   : in  std_logic_vector (31 downto 0);
    CLK : in  std_logic;
    Q   : out std_logic_vector (31 downto 0));
end entity fsqrt;

architecture rtl of fsqrt is

  function table(index: std_logic_vector(9 downto 0))
    return std_logic_vector
  is
    variable r : std_logic_vector(45 downto 0);
  begin
    case conv_integer(index) is
      when    0 => r := "1111111111000000000011100000000000111111111101";
      when    1 => r := "1111111101000000011011100000000010111111110101";
      when    2 => r := "1111111011000001001011100000000100111111100101";
      when    3 => r := "1111111001000010010011000000000110111111001101";
      when    4 => r := "1111110111000011110010000000001000111110101101";
      when    5 => r := "1111110101000101101000100000001010111110000101";
      when    6 => r := "1111110011000111110110100000001100111101010110";
      when    7 => r := "1111110001001010011011100000001110111100011110";
      when    8 => r := "1111101111001101011000000000010000111011011111";
      when    9 => r := "1111101101010000101011000000010010111010011000";
      when   10 => r := "1111101011010100010101100000010100111001001001";
      when   11 => r := "1111101001011000010110100000010110110111110011";
      when   12 => r := "1111100111011100101110100000011000110110010100";
      when   13 => r := "1111100101100001011100100000011010110100101110";
      when   14 => r := "1111100011100110100001100000011100110011000001";
      when   15 => r := "1111100001101011111101000000011110110001001011";
      when   16 => r := "1111011111110001101110100000100000101111001110";
      when   17 => r := "1111011101110111110110000000100010101101001001";
      when   18 => r := "1111011011111110010100000000100100101010111101";
      when   19 => r := "1111011010000101000111100000100110101000101001";
      when   20 => r := "1111011000001100010001000000101000100110001110";
      when   21 => r := "1111010110010011110000100000101010100011101011";
      when   22 => r := "1111010100011011100101100000101100100001000000";
      when   23 => r := "1111010010100011110000000000101110011110001110";
      when   24 => r := "1111010000101100010000000000110000011011010101";
      when   25 => r := "1111001110110101000101100000110010011000010011";
      when   26 => r := "1111001100111110010000000000110100010101001011";
      when   27 => r := "1111001011000111101111100000110110010001111100";
      when   28 => r := "1111001001010001100100100000111000001110100100";
      when   29 => r := "1111000111011011101110000000111010001011000110";
      when   30 => r := "1111000101100110001101000000111100000111100000";
      when   31 => r := "1111000011110001000000100000111110000011110010";
      when   32 => r := "1111000001111100001000100000111111111111111110";
      when   33 => r := "1111000000000111100101000001000001111100000010";
      when   34 => r := "1110111110010011010110000001000011110111111111";
      when   35 => r := "1110111100011111011011100001000101110011110101";
      when   36 => r := "1110111010101011110101100001000111101111100011";
      when   37 => r := "1110111000111000100011100001001001101011001010";
      when   38 => r := "1110110111000101100101100001001011100110101010";
      when   39 => r := "1110110101010010111100000001001101100010000010";
      when   40 => r := "1110110011100000100110000001001111011101010100";
      when   41 => r := "1110110001101110100100000001010001011000011111";
      when   42 => r := "1110101111111100110101100001010011010011100010";
      when   43 => r := "1110101110001011011011000001010101001110011110";
      when   44 => r := "1110101100011010010100000001010111001001010011";
      when   45 => r := "1110101010101001100000100001011001000100000001";
      when   46 => r := "1110101000111001000000000001011010111110101001";
      when   47 => r := "1110100111001000110011000001011100111001001001";
      when   48 => r := "1110100101011000111001100001011110110011100010";
      when   49 => r := "1110100011101001010011000001100000101101110100";
      when   50 => r := "1110100001111001111111100001100010100111111111";
      when   51 => r := "1110100000001010111111000001100100100010000011";
      when   52 => r := "1110011110011100010001100001100110011100000000";
      when   53 => r := "1110011100101101110110100001101000010101110111";
      when   54 => r := "1110011010111111101110100001101010001111100110";
      when   55 => r := "1110011001010001111001000001101100001001001111";
      when   56 => r := "1110010111100100010110100001101110000010110000";
      when   57 => r := "1110010101110111000110000001101111111100001011";
      when   58 => r := "1110010100001010001000000001110001110101011111";
      when   59 => r := "1110010010011101011100000001110011101110101101";
      when   60 => r := "1110010000110001000010100001110101100111110011";
      when   61 => r := "1110001111000100111011100001110111100000110010";
      when   62 => r := "1110001101011001000110000001111001011001101100";
      when   63 => r := "1110001011101101100011000001111011010010011110";
      when   64 => r := "1110001010000010010001100001111101001011001001";
      when   65 => r := "1110001000010111010010000001111111000011101110";
      when   66 => r := "1110000110101100100100100010000000111100001100";
      when   67 => r := "1110000101000010001000100010000010110100100011";
      when   68 => r := "1110000011010111111110000010000100101100110100";
      when   69 => r := "1110000001101110000101000010000110100100111110";
      when   70 => r := "1110000000000100011101100010001000011101000010";
      when   71 => r := "1101111110011011000111100010001010010100111111";
      when   72 => r := "1101111100110010000010100010001100001100110110";
      when   73 => r := "1101111011001001001111000010001110000100100110";
      when   74 => r := "1101111001100000101101000010001111111100001111";
      when   75 => r := "1101110111111000011011100010010001110011110010";
      when   76 => r := "1101110110010000011011100010010011101011001110";
      when   77 => r := "1101110100101000101100000010010101100010100100";
      when   78 => r := "1101110011000001001101100010010111011001110011";
      when   79 => r := "1101110001011010000000000010011001010000111100";
      when   80 => r := "1101101111110011000011000010011011000111111110";
      when   81 => r := "1101101110001100010111000010011100111110111010";
      when   82 => r := "1101101100100101111011000010011110110101110000";
      when   83 => r := "1101101010111111110000000010100000101100011111";
      when   84 => r := "1101101001011001110101100010100010100011001000";
      when   85 => r := "1101100111110100001011000010100100011001101010";
      when   86 => r := "1101100110001110110001000010100110010000000110";
      when   87 => r := "1101100100101001100111100010101000000110011100";
      when   88 => r := "1101100011000100101110000010101001111100101011";
      when   89 => r := "1101100001100000000100100010101011110010110100";
      when   90 => r := "1101011111111011101011000010101101101000110111";
      when   91 => r := "1101011110010111100001100010101111011110110100";
      when   92 => r := "1101011100110011101000000010110001010100101010";
      when   93 => r := "1101011011001111111110100010110011001010011010";
      when   94 => r := "1101011001101100100100100010110101000000000100";
      when   95 => r := "1101011000001001011010100010110110110101101000";
      when   96 => r := "1101010110100110011111100010111000101011000110";
      when   97 => r := "1101010101000011110101000010111010100000011101";
      when   98 => r := "1101010011100001011001100010111100010101101110";
      when   99 => r := "1101010001111111001101100010111110001010111001";
      when  100 => r := "1101010000011101010001000010111111111111111110";
      when  101 => r := "1101001110111011100011100011000001110100111101";
      when  102 => r := "1101001101011010000101100011000011101001110110";
      when  103 => r := "1101001011111000110111000011000101011110101000";
      when  104 => r := "1101001010010111110111100011000111010011010100";
      when  105 => r := "1101001000110111000111000011001001000111111011";
      when  106 => r := "1101000111010110100101100011001010111100011011";
      when  107 => r := "1101000101110110010010100011001100110000110110";
      when  108 => r := "1101000100010110001111000011001110100101001010";
      when  109 => r := "1101000010110110011010100011010000011001011000";
      when  110 => r := "1101000001010110110100100011010010001101100001";
      when  111 => r := "1100111111110111011101000011010100000001100100";
      when  112 => r := "1100111110011000010100100011010101110101100000";
      when  113 => r := "1100111100111001011010100011010111101001010110";
      when  114 => r := "1100111011011010101111000011011001011101000111";
      when  115 => r := "1100111001111100010010000011011011010000110010";
      when  116 => r := "1100111000011110000011100011011101000100010111";
      when  117 => r := "1100110111000000000011100011011110110111110101";
      when  118 => r := "1100110101100010010001100011100000101011001111";
      when  119 => r := "1100110100000100101110000011100010011110100010";
      when  120 => r := "1100110010100111011000100011100100010001101111";
      when  121 => r := "1100110001001010010001100011100110000100110111";
      when  122 => r := "1100101111101101011000000011100111110111111001";
      when  123 => r := "1100101110010000101101000011101001101010110101";
      when  124 => r := "1100101100110100010000000011101011011101101011";
      when  125 => r := "1100101011011000000001000011101101010000011011";
      when  126 => r := "1100101001111011111111100011101111000011000110";
      when  127 => r := "1100101000100000001100000011110000110101101011";
      when  128 => r := "1100100111000100100110100011110010101000001001";
      when  129 => r := "1100100101101001001110100011110100011010100011";
      when  130 => r := "1100100100001110000100000011110110001100110111";
      when  131 => r := "1100100010110011000111000011110111111111000101";
      when  132 => r := "1100100001011000011000000011111001110001001101";
      when  133 => r := "1100011111111101110110100011111011100011010000";
      when  134 => r := "1100011110100011100010000011111101010101001101";
      when  135 => r := "1100011101001001011011000011111111000111000101";
      when  136 => r := "1100011011101111100001100100000000111000110110";
      when  137 => r := "1100011010010101110101100100000010101010100010";
      when  138 => r := "1100011000111100010110100100000100011100001001";
      when  139 => r := "1100010111100011000100100100000110001101101010";
      when  140 => r := "1100010110001010000000000100000111111111000101";
      when  141 => r := "1100010100110001001000100100001001110000011011";
      when  142 => r := "1100010011011000011110000100001011100001101011";
      when  143 => r := "1100010010000000000000100100001101010010110110";
      when  144 => r := "1100010000100111110000000100001111000011111011";
      when  145 => r := "1100001111001111101100000100010000110100111011";
      when  146 => r := "1100001101110111110101100100010010100101110101";
      when  147 => r := "1100001100100000001011100100010100010110101010";
      when  148 => r := "1100001011001000101110000100010110000111011001";
      when  149 => r := "1100001001110001011101100100010111111000000011";
      when  150 => r := "1100001000011010011001100100011001101000101000";
      when  151 => r := "1100000111000011100010000100011011011001000111";
      when  152 => r := "1100000101101100110111000100011101001001100000";
      when  153 => r := "1100000100010110011001000100011110111001110100";
      when  154 => r := "1100000011000000000111000100100000101010000011";
      when  155 => r := "1100000001101010000001100100100010011010001100";
      when  156 => r := "1100000000010100001000100100100100001010010000";
      when  157 => r := "1011111110111110011100000100100101111010001111";
      when  158 => r := "1011111101101000111011100100100111101010001000";
      when  159 => r := "1011111100010011100111000100101001011001111100";
      when  160 => r := "1011111010111110011111000100101011001001101011";
      when  161 => r := "1011111001101001100011000100101100111001010100";
      when  162 => r := "1011111000010100110011100100101110101000110111";
      when  163 => r := "1011110111000000001111100100110000011000010110";
      when  164 => r := "1011110101101011111000000100110010000111101111";
      when  165 => r := "1011110100010111101100000100110011110111000100";
      when  166 => r := "1011110011000011101100000100110101100110010011";
      when  167 => r := "1011110001101111111000000100110111010101011100";
      when  168 => r := "1011110000011100010000000100111001000100100001";
      when  169 => r := "1011101111001000110011100100111010110011100000";
      when  170 => r := "1011101101110101100011000100111100100010011010";
      when  171 => r := "1011101100100010011110000100111110010001001110";
      when  172 => r := "1011101011001111100100100100111111111111111110";
      when  173 => r := "1011101001111100110111000101000001101110101000";
      when  174 => r := "1011101000101010010100100101000011011101001110";
      when  175 => r := "1011100111010111111110000101000101001011101110";
      when  176 => r := "1011100110000101110011000101000110111010001001";
      when  177 => r := "1011100100110011110011100101001000101000011110";
      when  178 => r := "1011100011100001111111000101001010010110101111";
      when  179 => r := "1011100010010000010110000101001100000100111011";
      when  180 => r := "1011100000111110111000100101001101110011000001";
      when  181 => r := "1011011111101101100110100101001111100001000010";
      when  182 => r := "1011011110011100011111000101010001001110111111";
      when  183 => r := "1011011101001011100011100101010010111100110110";
      when  184 => r := "1011011011111010110010100101010100101010101001";
      when  185 => r := "1011011010101010001101000101010110011000010110";
      when  186 => r := "1011011001011001110010100101011000000101111110";
      when  187 => r := "1011011000001001100011000101011001110011100001";
      when  188 => r := "1011010110111001011110100101011011100000111111";
      when  189 => r := "1011010101101001100101000101011101001110011000";
      when  190 => r := "1011010100011001110110100101011110111011101100";
      when  191 => r := "1011010011001010010011000101100000101000111011";
      when  192 => r := "1011010001111010111010000101100010010110000101";
      when  193 => r := "1011010000101011101100000101100100000011001011";
      when  194 => r := "1011001111011100101001000101100101110000001010";
      when  195 => r := "1011001110001101110000000101100111011101000110";
      when  196 => r := "1011001100111111000010100101101001001001111100";
      when  197 => r := "1011001011110000011111000101101010110110101110";
      when  198 => r := "1011001010100010000110100101101100100011011011";
      when  199 => r := "1011001001010011111000100101101110010000000010";
      when  200 => r := "1011001000000101110101000101101111111100100101";
      when  201 => r := "1011000110110111111100000101110001101001000011";
      when  202 => r := "1011000101101010001101100101110011010101011100";
      when  203 => r := "1011000100011100101001100101110101000001110000";
      when  204 => r := "1011000011001111010000000101110110101110000000";
      when  205 => r := "1011000010000010000000100101111000011010001010";
      when  206 => r := "1011000000110100111011100101111010000110010000";
      when  207 => r := "1010111111101000000001000101111011110010010001";
      when  208 => r := "1010111110011011010000100101111101011110001101";
      when  209 => r := "1010111101001110101010100101111111001010000100";
      when  210 => r := "1010111100000010001110100110000000110101110111";
      when  211 => r := "1010111010110101111100100110000010100001100100";
      when  212 => r := "1010111001101001110100100110000100001101001110";
      when  213 => r := "1010111000011101110111000110000101111000110010";
      when  214 => r := "1010110111010010000011100110000111100100010010";
      when  215 => r := "1010110110000110011001100110001001001111101101";
      when  216 => r := "1010110100111010111010000110001010111011000011";
      when  217 => r := "1010110011101111100100100110001100100110010100";
      when  218 => r := "1010110010100100011000100110001110010001100000";
      when  219 => r := "1010110001011001010110100110001111111100101000";
      when  220 => r := "1010110000001110011110100110010001100111101100";
      when  221 => r := "1010101111000011110000000110010011010010101010";
      when  222 => r := "1010101101111001001011100110010100111101100100";
      when  223 => r := "1010101100101110110000100110010110101000011010";
      when  224 => r := "1010101011100100011111100110011000010011001010";
      when  225 => r := "1010101010011010011000000110011001111101110110";
      when  226 => r := "1010101001010000011010100110011011101000011101";
      when  227 => r := "1010101000000110100110000110011101010011000000";
      when  228 => r := "1010100110111100111011100110011110111101011110";
      when  229 => r := "1010100101110011011010100110100000100111111000";
      when  230 => r := "1010100100101010000011000110100010010010001100";
      when  231 => r := "1010100011100000110100100110100011111100011101";
      when  232 => r := "1010100010010111110000000110100101100110101001";
      when  233 => r := "1010100001001110110101000110100111010000110000";
      when  234 => r := "1010100000000110000011000110101000111010110010";
      when  235 => r := "1010011110111101011010100110101010100100110001";
      when  236 => r := "1010011101110100111011000110101100001110101011";
      when  237 => r := "1010011100101100100101100110101101111000011111";
      when  238 => r := "1010011011100100011000100110101111100010010000";
      when  239 => r := "1010011010011100010101000110110001001011111100";
      when  240 => r := "1010011001010100011011000110110010110101100011";
      when  241 => r := "1010011000001100101010000110110100011111000110";
      when  242 => r := "1010010111000101000010000110110110001000100101";
      when  243 => r := "1010010101111101100011000110110111110001111111";
      when  244 => r := "1010010100110110001101100110111001011011010101";
      when  245 => r := "1010010011101111000000100110111011000100100110";
      when  246 => r := "1010010010100111111101000110111100101101110011";
      when  247 => r := "1010010001100001000010100110111110010110111011";
      when  248 => r := "1010010000011010010000100110111111111111111111";
      when  249 => r := "1010001111010011100111100111000001101000111110";
      when  250 => r := "1010001110001101001000000111000011010001111001";
      when  251 => r := "1010001101000110110000100111000100111010110000";
      when  252 => r := "1010001100000000100010100111000110100011100010";
      when  253 => r := "1010001010111010011101000111001000001100010000";
      when  254 => r := "1010001001110100100000100111001001110100111001";
      when  255 => r := "1010001000101110101100100111001011011101011110";
      when  256 => r := "1010000111101001000001100111001101000101111111";
      when  257 => r := "1010000110100011011111000111001110101110011011";
      when  258 => r := "1010000101011110000101000111010000010110110100";
      when  259 => r := "1010000100011000110100000111010001111111000111";
      when  260 => r := "1010000011010011101011100111010011100111010111";
      when  261 => r := "1010000010001110101011100111010101001111100010";
      when  262 => r := "1010000001001001110100000111010110110111101001";
      when  263 => r := "1010000000000101000101000111011000011111101011";
      when  264 => r := "1001111111000000011110100111011010000111101010";
      when  265 => r := "1001111101111100000001000111011011101111100011";
      when  266 => r := "1001111100110111101011100111011101010111011001";
      when  267 => r := "1001111011110011011110100111011110111111001010";
      when  268 => r := "1001111010101111011001100111100000100110110111";
      when  269 => r := "1001111001101011011101100111100010001110100000";
      when  270 => r := "1001111000100111101001100111100011110110000100";
      when  271 => r := "1001110111100011111110000111100101011101100101";
      when  272 => r := "1001110110100000011010100111100111000101000001";
      when  273 => r := "1001110101011100111111100111101000101100011001";
      when  274 => r := "1001110100011001101100100111101010010011101101";
      when  275 => r := "1001110011010110100010000111101011111010111100";
      when  276 => r := "1001110010010011011111100111101101100010000111";
      when  277 => r := "1001110001010000100101000111101111001001001111";
      when  278 => r := "1001110000001101110011000111110000110000010001";
      when  279 => r := "1001101111001011001000100111110010010111010001";
      when  280 => r := "1001101110001000100110100111110011111110001011";
      when  281 => r := "1001101101000110001100100111110101100101000010";
      when  282 => r := "1001101100000011111011000111110111001011110011";
      when  283 => r := "1001101011000001110001000111111000110010100010";
      when  284 => r := "1001101001111111101111000111111010011001001100";
      when  285 => r := "1001101000111101110101000111111011111111110010";
      when  286 => r := "1001100111111100000011000111111101100110010011";
      when  287 => r := "1001100110111010011000100111111111001100110010";
      when  288 => r := "1001100101111000110110101000000000110011001011";
      when  289 => r := "1001100100110111011100001000000010011001100000";
      when  290 => r := "1001100011110110001001001000000011111111110010";
      when  291 => r := "1001100010110100111110101000000101100101111111";
      when  292 => r := "1001100001110011111011101000000111001100001000";
      when  293 => r := "1001100000110011000000001000001000110010001110";
      when  294 => r := "1001011111110010001100101000001010011000001111";
      when  295 => r := "1001011110110001100000101000001011111110001100";
      when  296 => r := "1001011101110000111100101000001101100100000101";
      when  297 => r := "1001011100110000100000001000001111001001111010";
      when  298 => r := "1001011011110000001011001000010000101111101011";
      when  299 => r := "1001011010101111111110001000010010010101011000";
      when  300 => r := "1001011001101111111000001000010011111011000010";
      when  301 => r := "1001011000101111111010001000010101100000100110";
      when  302 => r := "1001010111110000000011101000010111000110000111";
      when  303 => r := "1001010110110000010100101000011000101011100100";
      when  304 => r := "1001010101110000101101001000011010010000111101";
      when  305 => r := "1001010100110001001101001000011011110110010010";
      when  306 => r := "1001010011110001110100001000011101011011100100";
      when  307 => r := "1001010010110010100011001000011111000000110001";
      when  308 => r := "1001010001110011011001001000100000100101111010";
      when  309 => r := "1001010000110100010111001000100010001010111111";
      when  310 => r := "1001001111110101011011101000100011110000000001";
      when  311 => r := "1001001110110110101000001000100101010100111110";
      when  312 => r := "1001001101110111111011101000100110111001110111";
      when  313 => r := "1001001100111001010110101000101000011110101101";
      when  314 => r := "1001001011111010111000101000101010000011011111";
      when  315 => r := "1001001010111100100010001000101011101000001100";
      when  316 => r := "1001001001111110010010101000101101001100110110";
      when  317 => r := "1001001001000000001010101000101110110001011100";
      when  318 => r := "1001001000000010001001101000110000010101111110";
      when  319 => r := "1001000111000100010000001000110001111010011100";
      when  320 => r := "1001000110000110011101001000110011011110110111";
      when  321 => r := "1001000101001000110001101000110101000011001101";
      when  322 => r := "1001000100001011001101001000110110100111100000";
      when  323 => r := "1001000011001101101111101000111000001011101111";
      when  324 => r := "1001000010010000011001101000111001101111111001";
      when  325 => r := "1001000001010011001010001000111011010100000001";
      when  326 => r := "1001000000010110000010001000111100111000000011";
      when  327 => r := "1000111111011001000000101000111110011100000011";
      when  328 => r := "1000111110011100000110101000111111111111111110";
      when  329 => r := "1000111101011111010011001001000001100011110111";
      when  330 => r := "1000111100100010100110101001000011000111101011";
      when  331 => r := "1000111011100110000001001001000100101011011011";
      when  332 => r := "1000111010101001100010101001000110001111000111";
      when  333 => r := "1000111001101101001010101001000111110010110000";
      when  334 => r := "1000111000110000111001101001001001010110010101";
      when  335 => r := "1000110111110100101111101001001010111001110110";
      when  336 => r := "1000110110111000101100101001001100011101010011";
      when  337 => r := "1000110101111100110000001001001110000000101101";
      when  338 => r := "1000110101000000111010001001001111100100000100";
      when  339 => r := "1000110100000101001011001001010001000111010110";
      when  340 => r := "1000110011001001100011001001010010101010100100";
      when  341 => r := "1000110010001110000001101001010100001101101111";
      when  342 => r := "1000110001010010100110101001010101110000110110";
      when  343 => r := "1000110000010111010010101001010111010011111001";
      when  344 => r := "1000101111011100000101001001011000110110111000";
      when  345 => r := "1000101110100000111110001001011010011001110100";
      when  346 => r := "1000101101100101111101101001011011111100101101";
      when  347 => r := "1000101100101011000100001001011101011111100001";
      when  348 => r := "1000101011110000010001001001011111000010010010";
      when  349 => r := "1000101010110101100100101001100000100100111111";
      when  350 => r := "1000101001111010111110101001100010000111101000";
      when  351 => r := "1000101001000000011111001001100011101010001110";
      when  352 => r := "1000101000000110000110001001100101001100110001";
      when  353 => r := "1000100111001011110011001001100110101111010000";
      when  354 => r := "1000100110010001100111001001101000010001101011";
      when  355 => r := "1000100101010111100001101001101001110100000010";
      when  356 => r := "1000100100011101100010101001101011010110010101";
      when  357 => r := "1000100011100011101001101001101100111000100101";
      when  358 => r := "1000100010101001110111001001101110011010110010";
      when  359 => r := "1000100001110000001011001001101111111100111011";
      when  360 => r := "1000100000110110100101101001110001011111000000";
      when  361 => r := "1000011111111101000110001001110011000001000001";
      when  362 => r := "1000011111000011101101001001110100100010111111";
      when  363 => r := "1000011110001010011010001001110110000100111010";
      when  364 => r := "1000011101010001001101101001110111100110110001";
      when  365 => r := "1000011100011000000111101001111001001000100100";
      when  366 => r := "1000011011011111000111101001111010101010010100";
      when  367 => r := "1000011010100110001101101001111100001100000000";
      when  368 => r := "1000011001101101011010001001111101101101101001";
      when  369 => r := "1000011000110100101101001001111111001111001101";
      when  370 => r := "1000010111111100000101101010000000110000101111";
      when  371 => r := "1000010111000011100100101010000010010010001101";
      when  372 => r := "1000010110001011001001101010000011110011101000";
      when  373 => r := "1000010101010010110101001010000101010100111110";
      when  374 => r := "1000010100011010100110001010000110110110010010";
      when  375 => r := "1000010011100010011101101010001000010111100010";
      when  376 => r := "1000010010101010011011001010001001111000101110";
      when  377 => r := "1000010001110010011110101010001011011001110111";
      when  378 => r := "1000010000111010101000001010001100111010111101";
      when  379 => r := "1000010000000010110111101010001110011011111111";
      when  380 => r := "1000001111001011001101001010001111111100111101";
      when  381 => r := "1000001110010011101000101010010001011101111000";
      when  382 => r := "1000001101011100001010001010010010111110110000";
      when  383 => r := "1000001100100100110001101010010100011111100100";
      when  384 => r := "1000001011101101011111001010010110000000010100";
      when  385 => r := "1000001010110110010010101010010111100001000001";
      when  386 => r := "1000001001111111001011101010011001000001101011";
      when  387 => r := "1000001001001000001010101010011010100010010001";
      when  388 => r := "1000001000010001001111101010011100000010110100";
      when  389 => r := "1000000111011010011010101010011101100011010011";
      when  390 => r := "1000000110100011101011001010011111000011101111";
      when  391 => r := "1000000101101101000001101010100000100100001000";
      when  392 => r := "1000000100110110011101101010100010000100011101";
      when  393 => r := "1000000100000000000000001010100011100100101110";
      when  394 => r := "1000000011001001100111101010100101000100111101";
      when  395 => r := "1000000010010011010101001010100110100101001000";
      when  396 => r := "1000000001011101001000101010101000000101001111";
      when  397 => r := "1000000000100111000001101010101001100101010011";
      when  398 => r := "0111111111110001000000001010101011000101010100";
      when  399 => r := "0111111110111011000100101010101100100101010010";
      when  400 => r := "0111111110000101001110101010101110000101001100";
      when  401 => r := "0111111101001111011110101010101111100101000010";
      when  402 => r := "0111111100011001110100001010110001000100110101";
      when  403 => r := "0111111011100100001111001010110010100100100101";
      when  404 => r := "0111111010101110101111101010110100000100010010";
      when  405 => r := "0111111001111001010110001010110101100011111011";
      when  406 => r := "0111111001000100000001101010110111000011100001";
      when  407 => r := "0111111000001110110011001010111000100011000100";
      when  408 => r := "0111110111011001101010001010111010000010100011";
      when  409 => r := "0111110110100100100110101010111011100001111111";
      when  410 => r := "0111110101101111101000101010111101000001010111";
      when  411 => r := "0111110100111010110000001010111110100000101101";
      when  412 => r := "0111110100000101111101001010111111111111111111";
      when  413 => r := "0111110011010001001111101011000001011111001110";
      when  414 => r := "0111110010011100100111101011000010111110011001";
      when  415 => r := "0111110001101000000101001011000100011101100001";
      when  416 => r := "0111110000110011100111101011000101111100100110";
      when  417 => r := "0111101111111111010000001011000111011011100111";
      when  418 => r := "0111101111001010111101101011001000111010100110";
      when  419 => r := "0111101110010110110000101011001010011001100001";
      when  420 => r := "0111101101100010101001001011001011111000011001";
      when  421 => r := "0111101100101110100111001011001101010111001101";
      when  422 => r := "0111101011111010101010001011001110110101111111";
      when  423 => r := "0111101011000110110010101011010000010100101101";
      when  424 => r := "0111101010010011000000001011010001110011011000";
      when  425 => r := "0111101001011111010011101011010011010001111111";
      when  426 => r := "0111101000101011101011101011010100110000100100";
      when  427 => r := "0111100111111000001001101011010110001111000100";
      when  428 => r := "0111100111000100101100001011010111101101100011";
      when  429 => r := "0111100110010001010100101011011001001011111101";
      when  430 => r := "0111100101011110000010001011011010101010010100";
      when  431 => r := "0111100100101010110100101011011100001000101001";
      when  432 => r := "0111100011110111101100001011011101100110111010";
      when  433 => r := "0111100011000100101001001011011111000101001000";
      when  434 => r := "0111100010010001101011101011100000100011010010";
      when  435 => r := "0111100001011110110011001011100010000001011010";
      when  436 => r := "0111100000101011111111101011100011011111011110";
      when  437 => r := "0111011111111001010001001011100100111101011111";
      when  438 => r := "0111011111000110100111101011100110011011011110";
      when  439 => r := "0111011110010100000011101011100111111001011001";
      when  440 => r := "0111011101100001100100101011101001010111010000";
      when  441 => r := "0111011100101111001010101011101010110101000101";
      when  442 => r := "0111011011111100110110001011101100010010110110";
      when  443 => r := "0111011011001010100110001011101101110000100100";
      when  444 => r := "0111011010011000011011001011101111001110010000";
      when  445 => r := "0111011001100110010101101011110000101011110111";
      when  446 => r := "0111011000110100010101001011110010001001011100";
      when  447 => r := "0111011000000010011001001011110011100110111110";
      when  448 => r := "0111010111010000100010101011110101000100011100";
      when  449 => r := "0111010110011110110000101011110110100001111000";
      when  450 => r := "0111010101101101000100001011110111111111010000";
      when  451 => r := "0111010100111011011100001011111001011100100101";
      when  452 => r := "0111010100001001111001001011111010111001111000";
      when  453 => r := "0111010011011000011011001011111100010111000111";
      when  454 => r := "0111010010100111000010001011111101110100010011";
      when  455 => r := "0111010001110101101110001011111111010001011100";
      when  456 => r := "0111010001000100011111001100000000101110100001";
      when  457 => r := "0111010000010011010100101100000010001011100100";
      when  458 => r := "0111001111100010001111001100000011101000100100";
      when  459 => r := "0111001110110001001110001100000101000101100001";
      when  460 => r := "0111001110000000010010101100000110100010011010";
      when  461 => r := "0111001101001111011011101100000111111111010000";
      when  462 => r := "0111001100011110101001101100001001011100000011";
      when  463 => r := "0111001011101101111100001100001010111000110100";
      when  464 => r := "0111001010111101010011101100001100010101100001";
      when  465 => r := "0111001010001100101111101100001101110010001100";
      when  466 => r := "0111001001011100010000101100001111001110110011";
      when  467 => r := "0111001000101011110110001100010000101011011000";
      when  468 => r := "0111000111111011100000101100010010000111111001";
      when  469 => r := "0111000111001011010000001100010011100100010111";
      when  470 => r := "0111000110011011000100001100010101000000110010";
      when  471 => r := "0111000101101010111100101100010110011101001010";
      when  472 => r := "0111000100111010111001101100010111111001100000";
      when  473 => r := "0111000100001010111011101100011001010101110010";
      when  474 => r := "0111000011011011000010101100011010110010000001";
      when  475 => r := "0111000010101011001101101100011100001110001101";
      when  476 => r := "0111000001111011011101101100011101101010010110";
      when  477 => r := "0111000001001011110010001100011111000110011101";
      when  478 => r := "0111000000011100001011101100100000100010100000";
      when  479 => r := "0110111111101100101001001100100001111110100000";
      when  480 => r := "0110111110111101001011101100100011011010011110";
      when  481 => r := "0110111110001101110010101100100100110110011000";
      when  482 => r := "0110111101011110011110001100100110010010010000";
      when  483 => r := "0110111100101111001110101100100111101110000011";
      when  484 => r := "0110111100000000000011001100101001001001110101";
      when  485 => r := "0110111011010000111100101100101010100101100011";
      when  486 => r := "0110111010100001111010001100101100000001001111";
      when  487 => r := "0110111001110010111100101100101101011100111000";
      when  488 => r := "0110111001000100000011001100101110111000011110";
      when  489 => r := "0110111000010101001110101100110000010100000000";
      when  490 => r := "0110110111100110011110001100110001101111100001";
      when  491 => r := "0110110110110111110010101100110011001010111101";
      when  492 => r := "0110110110001001001011001100110100100110011000";
      when  493 => r := "0110110101011010101000101100110110000001101110";
      when  494 => r := "0110110100101100001010001100110111011101000010";
      when  495 => r := "0110110011111101110000001100111000111000010100";
      when  496 => r := "0110110011001111011010101100111010010011100010";
      when  497 => r := "0110110010100001001001101100111011101110101101";
      when  498 => r := "0110110001110010111100101100111101001001110111";
      when  499 => r := "0110110001000100110100101100111110100100111100";
      when  500 => r := "0110110000010110110000101100111111111111111111";
      when  501 => r := "0110101111101000110000101101000001011010111111";
      when  502 => r := "0110101110111010110101101101000010110101111100";
      when  503 => r := "0110101110001100111110101101000100010000110110";
      when  504 => r := "0110101101011111001100001101000101101011101101";
      when  505 => r := "0110101100110001011101101101000111000110100010";
      when  506 => r := "0110101100000011110011101101001000100001010100";
      when  507 => r := "0110101011010110001110001101001001111100000011";
      when  508 => r := "0110101010101000101100101101001011010110101111";
      when  509 => r := "0110101001111011001111101101001100110001011000";
      when  510 => r := "0110101001001101110111001101001110001011111110";
      when  511 => r := "0110101000100000100010001101001111100110100010";
      when  512 => r := "0110100111011100101100001101010001101110001111";
      when  513 => r := "0110100110000010011100001101010100100011000110";
      when  514 => r := "0110100100101000011101101101010111010111110000";
      when  515 => r := "0110100011001110101111001101011010001100010000";
      when  516 => r := "0110100001110101010010001101011101000000100100";
      when  517 => r := "0110100000011100000101001101011111110100101101";
      when  518 => r := "0110011111000011001001001101100010101000101010";
      when  519 => r := "0110011101101010011101001101100101011100011110";
      when  520 => r := "0110011100010010000001101101101000010000000110";
      when  521 => r := "0110011010111001110110101101101011000011100010";
      when  522 => r := "0110011001100001111011101101101101110110110100";
      when  523 => r := "0110011000001010010000101101110000101001111011";
      when  524 => r := "0110010110110010110101101101110011011100110111";
      when  525 => r := "0110010101011011101011001101110110001111100111";
      when  526 => r := "0110010100000100110000001101111001000010001110";
      when  527 => r := "0110010010101110000101001101111011110100101001";
      when  528 => r := "0110010001010111101001101101111110100110111001";
      when  529 => r := "0110010000000001011110001110000001011000111111";
      when  530 => r := "0110001110101011100010001110000100001010111001";
      when  531 => r := "0110001101010101110101101110000110111100101001";
      when  532 => r := "0110001100000000011000101110001001101110001111";
      when  533 => r := "0110001010101011001010101110001100011111101010";
      when  534 => r := "0110001001010110001100001110001111010000111010";
      when  535 => r := "0110001000000001011101001110010010000001111111";
      when  536 => r := "0110000110101100111101001110010100110010111010";
      when  537 => r := "0110000101011000101100101110010111100011101010";
      when  538 => r := "0110000100000100101010101110011010010100010000";
      when  539 => r := "0110000010110000110111101110011101000100101100";
      when  540 => r := "0110000001011101010011101110011111110100111101";
      when  541 => r := "0110000000001001111110101110100010100101000011";
      when  542 => r := "0101111110110110111000001110100101010100111111";
      when  543 => r := "0101111101100100000000101110101000000100110000";
      when  544 => r := "0101111100010001010111001110101010110100011001";
      when  545 => r := "0101111010111110111100101110101101100011110110";
      when  546 => r := "0101111001101100110000101110110000010011001000";
      when  547 => r := "0101111000011010110011001110110011000010010000";
      when  548 => r := "0101110111001001000011101110110101110001001111";
      when  549 => r := "0101110101110111100010101110111000100000000011";
      when  550 => r := "0101110100100110010000001110111011001110101100";
      when  551 => r := "0101110011010101001011001110111101111101001101";
      when  552 => r := "0101110010000100010100101111000000101011100010";
      when  553 => r := "0101110000110011101100001111000011011001101110";
      when  554 => r := "0101101111100011010001101111000110000111101111";
      when  555 => r := "0101101110010011000101001111001000110101100110";
      when  556 => r := "0101101101000011000110001111001011100011010100";
      when  557 => r := "0101101011110011010101001111001110010000110111";
      when  558 => r := "0101101010100011110010001111010000111110010000";
      when  559 => r := "0101101001010100011100001111010011101011100000";
      when  560 => r := "0101101000000101010100001111010110011000100110";
      when  561 => r := "0101100110110110011001101111011001000101100010";
      when  562 => r := "0101100101100111101100101111011011110010010011";
      when  563 => r := "0101100100011001001101001111011110011110111011";
      when  564 => r := "0101100011001010111010101111100001001011011010";
      when  565 => r := "0101100001111100110101101111100011110111101110";
      when  566 => r := "0101100000101110111110001111100110100011111001";
      when  567 => r := "0101011111100001010011101111101001001111111001";
      when  568 => r := "0101011110010011110110001111101011111011110001";
      when  569 => r := "0101011101000110100101101111101110100111011111";
      when  570 => r := "0101011011111001100010001111110001010011000011";
      when  571 => r := "0101011010101100101100001111110011111110011101";
      when  572 => r := "0101011001100000000010101111110110101001101101";
      when  573 => r := "0101011000010011100101101111111001010100110101";
      when  574 => r := "0101010111000111010101101111111011111111110011";
      when  575 => r := "0101010101111011010010101111111110101010100111";
      when  576 => r := "0101010100101111011100010000000001010101010001";
      when  577 => r := "0101010011100011110010010000000011111111110011";
      when  578 => r := "0101010010011000010100110000000110101010001011";
      when  579 => r := "0101010001001101000100010000001001010100011000";
      when  580 => r := "0101010000000001111111110000001011111110011110";
      when  581 => r := "0101001110110111000111110000001110101000011001";
      when  582 => r := "0101001101101100011100010000010001010010001011";
      when  583 => r := "0101001100100001111100110000010011111011110100";
      when  584 => r := "0101001011010111101001110000010110100101010100";
      when  585 => r := "0101001010001101100010110000011001001110101010";
      when  586 => r := "0101001001000011100111110000011011110111111000";
      when  587 => r := "0101000111111001111001010000011110100000111011";
      when  588 => r := "0101000110110000010110010000100001001001110110";
      when  589 => r := "0101000101100110111111110000100011110010100111";
      when  590 => r := "0101000100011101110101010000100110011011001111";
      when  591 => r := "0101000011010100110110010000101001000011101111";
      when  592 => r := "0101000010001100000011010000101011101100000101";
      when  593 => r := "0101000001000011011011110000101110010100010010";
      when  594 => r := "0100111111111011000000010000110000111100010110";
      when  595 => r := "0100111110110010110000010000110011100100010001";
      when  596 => r := "0100111101101010101100010000110110001100000010";
      when  597 => r := "0100111100100010110011110000111000110011101011";
      when  598 => r := "0100111011011011000110010000111011011011001100";
      when  599 => r := "0100111010010011100100110000111110000010100010";
      when  600 => r := "0100111001001100001110110001000000101001110000";
      when  601 => r := "0100111000000101000011110001000011010000110101";
      when  602 => r := "0100110110111110000100010001000101110111110010";
      when  603 => r := "0100110101110111010000010001001000011110100101";
      when  604 => r := "0100110100110000100111010001001011000101001111";
      when  605 => r := "0100110011101010001001110001001101101011110001";
      when  606 => r := "0100110010100011110111010001010000010010001001";
      when  607 => r := "0100110001011101101111110001010010111000011010";
      when  608 => r := "0100110000010111110011010001010101011110100001";
      when  609 => r := "0100101111010010000001110001011000000100100000";
      when  610 => r := "0100101110001100011011110001011010101010010101";
      when  611 => r := "0100101101000111000000010001011101010000000011";
      when  612 => r := "0100101100000001101111110001011111110101100111";
      when  613 => r := "0100101010111100101001110001100010011011000100";
      when  614 => r := "0100101001110111101111010001100101000000010110";
      when  615 => r := "0100101000110010111110110001100111100101100010";
      when  616 => r := "0100100111101110011001010001101010001010100100";
      when  617 => r := "0100100110101001111110110001101100101111011101";
      when  618 => r := "0100100101100101101110110001101111010100001101";
      when  619 => r := "0100100100100001101000110001110001111000110111";
      when  620 => r := "0100100011011101101101110001110100011101010111";
      when  621 => r := "0100100010011001111101010001110111000001101110";
      when  622 => r := "0100100001010110010111010001111001100101111101";
      when  623 => r := "0100100000010010111011110001111100001010000011";
      when  624 => r := "0100011111001111101010010001111110101110000010";
      when  625 => r := "0100011110001100100011010010000001010001111000";
      when  626 => r := "0100011101001001100110110010000011110101100101";
      when  627 => r := "0100011100000110110100010010000110011001001010";
      when  628 => r := "0100011011000100001100010010001000111100100110";
      when  629 => r := "0100011010000001101101110010001011011111111011";
      when  630 => r := "0100011000111111011001110010001110000011000111";
      when  631 => r := "0100010111111101010000010010010000100110001010";
      when  632 => r := "0100010110111011010000010010010011001001000110";
      when  633 => r := "0100010101111001011010110010010101101011111001";
      when  634 => r := "0100010100110111101110110010011000001110100100";
      when  635 => r := "0100010011110110001100110010011010110001000111";
      when  636 => r := "0100010010110100110100110010011101010011100010";
      when  637 => r := "0100010001110011100110110010011111110101110100";
      when  638 => r := "0100010000110010100010010010100010010111111111";
      when  639 => r := "0100001111110001100111110010100100111010000001";
      when  640 => r := "0100001110110000110110110010100111011011111011";
      when  641 => r := "0100001101110000001111110010101001111101101101";
      when  642 => r := "0100001100101111110010010010101100011111010111";
      when  643 => r := "0100001011101111011110010010101111000000111001";
      when  644 => r := "0100001010101111010011110010110001100010010100";
      when  645 => r := "0100001001101111010011010010110100000011100101";
      when  646 => r := "0100001000101111011011110010110110100100101111";
      when  647 => r := "0100000111101111101110010010111001000101110001";
      when  648 => r := "0100000110110000001001110010111011100110101011";
      when  649 => r := "0100000101110000101110110010111110000111011101";
      when  650 => r := "0100000100110001011101010011000000101000000111";
      when  651 => r := "0100000011110010010100110011000011001000101010";
      when  652 => r := "0100000010110011010101110011000101101001000100";
      when  653 => r := "0100000001110100100000010011001000001001010110";
      when  654 => r := "0100000000110101110011110011001010101001100001";
      when  655 => r := "0011111111110111010000010011001101001001100100";
      when  656 => r := "0011111110111000110110010011001111101001011111";
      when  657 => r := "0011111101111010100101010011010010001001010010";
      when  658 => r := "0011111100111100011101010011010100101000111110";
      when  659 => r := "0011111011111110011110010011010111001000100010";
      when  660 => r := "0011111011000000101000110011011001100111111101";
      when  661 => r := "0011111010000010111011110011011100000111010001";
      when  662 => r := "0011111001000101010111110011011110100110011110";
      when  663 => r := "0011111000000111111100110011100001000101100010";
      when  664 => r := "0011110111001010101010010011100011100100100000";
      when  665 => r := "0011110110001101100001010011100110000011010101";
      when  666 => r := "0011110101010000100000110011101000100010000011";
      when  667 => r := "0011110100010011101000110011101011000000101010";
      when  668 => r := "0011110011010110111001110011101101011111001000";
      when  669 => r := "0011110010011010010011010011101111111101100000";
      when  670 => r := "0011110001011101110101110011110010011011101111";
      when  671 => r := "0011110000100001100000110011110100111001110111";
      when  672 => r := "0011101111100101010100110011110111010111110111";
      when  673 => r := "0011101110101001010000110011111001110101110000";
      when  674 => r := "0011101101101101010101110011111100010011100001";
      when  675 => r := "0011101100110001100010110011111110110001001100";
      when  676 => r := "0011101011110101111000110100000001001110101110";
      when  677 => r := "0011101010111010010110110100000011101100001001";
      when  678 => r := "0011101001111110111101110100000110001001011100";
      when  679 => r := "0011101001000011101100110100001000100110101000";
      when  680 => r := "0011101000001000100100010100001011000011101101";
      when  681 => r := "0011100111001101100011110100001101100000101011";
      when  682 => r := "0011100110010010101011110100001111111101100001";
      when  683 => r := "0011100101010111111100010100010010011010001111";
      when  684 => r := "0011100100011101010100110100010100110110110111";
      when  685 => r := "0011100011100010110101110100010111010011010110";
      when  686 => r := "0011100010101000011110110100011001101111101111";
      when  687 => r := "0011100001101110001111110100011100001100000001";
      when  688 => r := "0011100000110100001000110100011110101000001011";
      when  689 => r := "0011011111111010001010010100100001000100001110";
      when  690 => r := "0011011111000000010011110100100011100000001001";
      when  691 => r := "0011011110000110100101010100100101111011111110";
      when  692 => r := "0011011101001100111110110100101000010111101011";
      when  693 => r := "0011011100010011011111110100101010110011010010";
      when  694 => r := "0011011011011010001001010100101101001110110000";
      when  695 => r := "0011011010100000111010110100101111101010000111";
      when  696 => r := "0011011001100111110011110100110010000101011000";
      when  697 => r := "0011011000101110110100110100110100100000100010";
      when  698 => r := "0011010111110101111101110100110110111011100100";
      when  699 => r := "0011010110111101001110010100111001010110100000";
      when  700 => r := "0011010110000100100110110100111011110001010100";
      when  701 => r := "0011010101001100000111010100111110001100000000";
      when  702 => r := "0011010100010011101110110101000000100110100111";
      when  703 => r := "0011010011011011011110110101000011000001000101";
      when  704 => r := "0011010010100011010101110101000101011011011110";
      when  705 => r := "0011010001101011010100110101000111110101101110";
      when  706 => r := "0011010000110011011011010101001010001111111001";
      when  707 => r := "0011001111111011101001110101001100101001111010";
      when  708 => r := "0011001111000011111111010101001111000011110111";
      when  709 => r := "0011001110001100011100010101010001011101101101";
      when  710 => r := "0011001101010101000001010101010011110111011010";
      when  711 => r := "0011001100011101101101010101010110010001000010";
      when  712 => r := "0011001011100110100001010101011000101010100001";
      when  713 => r := "0011001010101111011100010101011011000011111011";
      when  714 => r := "0011001001111000011110110101011101011101001101";
      when  715 => r := "0011001001000001101000110101011111110110011001";
      when  716 => r := "0011001000001010111001110101100010001111011110";
      when  717 => r := "0011000111010100010010010101100100101000011100";
      when  718 => r := "0011000110011101110010010101100111000001010011";
      when  719 => r := "0011000101100111011001010101101001011010000100";
      when  720 => r := "0011000100110001000111110101101011110010101101";
      when  721 => r := "0011000011111010111101010101101110001011010000";
      when  722 => r := "0011000011000100111010010101110000100011101100";
      when  723 => r := "0011000010001110111110010101110010111100000001";
      when  724 => r := "0011000001011001001001010101110101010100010000";
      when  725 => r := "0011000000100011011011110101110111101100011000";
      when  726 => r := "0010111111101101110100110101111010000100011010";
      when  727 => r := "0010111110111000010101010101111100011100010100";
      when  728 => r := "0010111110000010111100110101111110110100001000";
      when  729 => r := "0010111101001101101011010110000001001011110101";
      when  730 => r := "0010111100011000100000110110000011100011011011";
      when  731 => r := "0010111011100011011101010110000101111010111011";
      when  732 => r := "0010111010101110100000110110001000010010010100";
      when  733 => r := "0010111001111001101011010110001010101001100110";
      when  734 => r := "0010111001000100111100110110001101000000110001";
      when  735 => r := "0010111000010000010100110110001111010111110111";
      when  736 => r := "0010110111011011110011110110010001101110110110";
      when  737 => r := "0010110110100111011001110110010100000101101110";
      when  738 => r := "0010110101110011000110010110010110011100100000";
      when  739 => r := "0010110100111110111001110110011000110011001011";
      when  740 => r := "0010110100001010110100010110011011001001101111";
      when  741 => r := "0010110011010110110101010110011101100000001101";
      when  742 => r := "0010110010100010111100110110011111110110100101";
      when  743 => r := "0010110001101111001011010110100010001100110110";
      when  744 => r := "0010110000111011100000010110100100100011000001";
      when  745 => r := "0010110000000111111100010110100110111001000101";
      when  746 => r := "0010101111010100011110010110101001001111000100";
      when  747 => r := "0010101110100001000111010110101011100100111011";
      when  748 => r := "0010101101101101110111010110101101111010101011";
      when  749 => r := "0010101100111010101101010110110000010000010110";
      when  750 => r := "0010101100000111101001110110110010100101111011";
      when  751 => r := "0010101011010100101101010110110100111011011000";
      when  752 => r := "0010101010100001110110110110110111010000110000";
      when  753 => r := "0010101001101111000111010110111001100110000000";
      when  754 => r := "0010101000111100011101110110111011111011001011";
      when  755 => r := "0010101000001001111010110110111110010000010000";
      when  756 => r := "0010100111010111011110010111000000100101001110";
      when  757 => r := "0010100110100101001000010111000010111010000110";
      when  758 => r := "0010100101110010111000110111000101001110110110";
      when  759 => r := "0010100101000000101111010111000111100011100010";
      when  760 => r := "0010100100001110101100010111001001111000000111";
      when  761 => r := "0010100011011100101111110111001100001100100101";
      when  762 => r := "0010100010101010111001010111001110100000111110";
      when  763 => r := "0010100001111001001000110111010000110101010001";
      when  764 => r := "0010100001000111011111010111010011001001011100";
      when  765 => r := "0010100000010101111011010111010101011101100011";
      when  766 => r := "0010011111100100011101110111010111110001100011";
      when  767 => r := "0010011110110011000110110111011010000101011011";
      when  768 => r := "0010011110000001110101110111011100011001001110";
      when  769 => r := "0010011101010000101010110111011110101100111011";
      when  770 => r := "0010011100011111100101110111100001000000100011";
      when  771 => r := "0010011011101110100111010111100011010100000011";
      when  772 => r := "0010011010111101101110010111100101100111011111";
      when  773 => r := "0010011010001100111011110111100111111010110100";
      when  774 => r := "0010011001011100001111010111101010001110000010";
      when  775 => r := "0010011000101011101000110111101100100001001011";
      when  776 => r := "0010010111111011001000010111101110110100001101";
      when  777 => r := "0010010111001010101101110111110001000111001010";
      when  778 => r := "0010010110011010011001010111110011011010000000";
      when  779 => r := "0010010101101010001010110111110101101100110000";
      when  780 => r := "0010010100111010000010010111110111111111011010";
      when  781 => r := "0010010100001001111111110111111010010001111110";
      when  782 => r := "0010010011011010000010110111111100100100011100";
      when  783 => r := "0010010010101010001011110111111110110110110101";
      when  784 => r := "0010010001111010011010111000000001001001000111";
      when  785 => r := "0010010001001010101111011000000011011011010100";
      when  786 => r := "0010010000011011001010011000000101101101011001";
      when  787 => r := "0010001111101011101010011000000111111111011011";
      when  788 => r := "0010001110111100010000111000001010010001010100";
      when  789 => r := "0010001110001100111100111000001100100011001001";
      when  790 => r := "0010001101011101101110011000001110110100111000";
      when  791 => r := "0010001100101110100101111000010001000110100000";
      when  792 => r := "0010001011111111100010111000010011011000000100";
      when  793 => r := "0010001011010000100101111000010101101001100000";
      when  794 => r := "0010001010100001101110011000010111111010110111";
      when  795 => r := "0010001001110010111100011000011010001100001001";
      when  796 => r := "0010001001000100010000011000011100011101010100";
      when  797 => r := "0010001000010101101001011000011110101110011011";
      when  798 => r := "0010000111100111001000111000100000111111011001";
      when  799 => r := "0010000110111000101101011000100011010000010011";
      when  800 => r := "0010000110001010010111011000100101100001001000";
      when  801 => r := "0010000101011100000111011000100111110001110110";
      when  802 => r := "0010000100101101111100011000101010000010011111";
      when  803 => r := "0010000011111111110111011000101100010011000001";
      when  804 => r := "0010000011010001110111011000101110100011011111";
      when  805 => r := "0010000010100011111101011000110000110011110110";
      when  806 => r := "0010000001110110001000011000110011000100001000";
      when  807 => r := "0010000001001000011001011000110101010100010011";
      when  808 => r := "0010000000011010101111011000110111100100011010";
      when  809 => r := "0001111111101101001010111000111001110100011010";
      when  810 => r := "0001111110111111101011111000111100000100010101";
      when  811 => r := "0001111110010010010001111000111110010100001011";
      when  812 => r := "0001111101100100111101111001000000100011111010";
      when  813 => r := "0001111100110111101110111001000010110011100011";
      when  814 => r := "0001111100001010100101011001000101000011000111";
      when  815 => r := "0001111011011101100000111001000111010010100110";
      when  816 => r := "0001111010110000100001111001001001100001111111";
      when  817 => r := "0001111010000011100111111001001011110001010011";
      when  818 => r := "0001111001010110110011011001001110000000100001";
      when  819 => r := "0001111000101010000100011001010000001111101000";
      when  820 => r := "0001110111111101011010011001010010011110101011";
      when  821 => r := "0001110111010000110101011001010100101101101000";
      when  822 => r := "0001110110100100010101111001010110111100100000";
      when  823 => r := "0001110101110111111011111001011001001011010000";
      when  824 => r := "0001110101001011100110011001011011011001111101";
      when  825 => r := "0001110100011111010110011001011101101000100100";
      when  826 => r := "0001110011110011001011011001011111110111000101";
      when  827 => r := "0001110011000111000101111001100010000101100000";
      when  828 => r := "0001110010011011000101011001100100010011110110";
      when  829 => r := "0001110001101111001001011001100110100010001000";
      when  830 => r := "0001110001000011010010111001101000110000010011";
      when  831 => r := "0001110000010111100001111001101010111110010111";
      when  832 => r := "0001101111101011110101011001101101001100011000";
      when  833 => r := "0001101111000000001101111001101111011010010011";
      when  834 => r := "0001101110010100101011011001110001101000001001";
      when  835 => r := "0001101101101001001110011001110011110101111000";
      when  836 => r := "0001101100111101110101111001110110000011100011";
      when  837 => r := "0001101100010010100010111001111000010001000111";
      when  838 => r := "0001101011100111010100011001111010011110100111";
      when  839 => r := "0001101010111100001010111001111100101100000001";
      when  840 => r := "0001101010010001000110011001111110111001010110";
      when  841 => r := "0001101001100110000110111010000001000110100101";
      when  842 => r := "0001101000111011001011111010000011010011110000";
      when  843 => r := "0001101000010000010110011010000101100000110100";
      when  844 => r := "0001100111100101100101011010000111101101110011";
      when  845 => r := "0001100110111010111000111010001001111010101111";
      when  846 => r := "0001100110010000010001111010001100000111100011";
      when  847 => r := "0001100101100101101111011010001110010100010010";
      when  848 => r := "0001100100111011010001111010010000100000111100";
      when  849 => r := "0001100100010000111000111010010010101101100001";
      when  850 => r := "0001100011100110100100111010010100111010000001";
      when  851 => r := "0001100010111100010101111010010111000110011010";
      when  852 => r := "0001100010010010001011011010011001010010101111";
      when  853 => r := "0001100001101000000101011010011011011111000000";
      when  854 => r := "0001100000111110000100011010011101101011001010";
      when  855 => r := "0001100000010100001000011010011111110111001110";
      when  856 => r := "0001011111101010010000011010100010000011001111";
      when  857 => r := "0001011111000000011101111010100100001111001001";
      when  858 => r := "0001011110010110101111011010100110011010111111";
      when  859 => r := "0001011101101101000101111010101000100110101111";
      when  860 => r := "0001011101000011100000111010101010110010011010";
      when  861 => r := "0001011100011010000000111010101100111101111111";
      when  862 => r := "0001011011110000100100111010101111001001100001";
      when  863 => r := "0001011011000111001101111010110001010100111100";
      when  864 => r := "0001011010011101111011011010110011100000010011";
      when  865 => r := "0001011001110100101101011010110101101011100100";
      when  866 => r := "0001011001001011100100011010110111110110101111";
      when  867 => r := "0001011000100010011111011010111010000001110111";
      when  868 => r := "0001010111111001011111011010111100001100111000";
      when  869 => r := "0001010111010000100011011010111110010111110101";
      when  870 => r := "0001010110100111101100011011000000100010101100";
      when  871 => r := "0001010101111110111001111011000010101101011110";
      when  872 => r := "0001010101010110001011011011000100111000001101";
      when  873 => r := "0001010100101101100001111011000111000010110100";
      when  874 => r := "0001010100000100111100011011001001001101011000";
      when  875 => r := "0001010011011100011011111011001011010111110101";
      when  876 => r := "0001010010110011111111011011001101100010001111";
      when  877 => r := "0001010010001011100111011011001111101100100011";
      when  878 => r := "0001010001100011010011111011010001110110110010";
      when  879 => r := "0001010000111011000100111011010100000000111011";
      when  880 => r := "0001010000010010111010011011010110001010111111";
      when  881 => r := "0001001111101010110011111011011000010101000000";
      when  882 => r := "0001001111000010110001111011011010011110111011";
      when  883 => r := "0001001110011010110100011011011100101000110000";
      when  884 => r := "0001001101110010111010111011011110110010100010";
      when  885 => r := "0001001101001011000101111011100000111100001110";
      when  886 => r := "0001001100100011010101011011100011000101110100";
      when  887 => r := "0001001011111011101000111011100101001111010110";
      when  888 => r := "0001001011010100000000111011100111011000110011";
      when  889 => r := "0001001010101100011100111011101001100010001100";
      when  890 => r := "0001001010000100111101011011101011101011011111";
      when  891 => r := "0001001001011101100010011011101101110100101100";
      when  892 => r := "0001001000110110001011011011101111111101110101";
      when  893 => r := "0001001000001110111000011011110010000110111010";
      when  894 => r := "0001000111100111101001111011110100001111111001";
      when  895 => r := "0001000111000000011111011011110110011000110100";
      when  896 => r := "0001000110011001011001011011111000100001101001";
      when  897 => r := "0001000101110010010111011011111010101010011010";
      when  898 => r := "0001000101001011011001011011111100110011000111";
      when  899 => r := "0001000100100100011111111011111110111011101101";
      when  900 => r := "0001000011111101101010011100000001000100001111";
      when  901 => r := "0001000011010110111000111100000011001100101101";
      when  902 => r := "0001000010110000001011111100000101010101000100";
      when  903 => r := "0001000010001001100010011100000111011101011001";
      when  904 => r := "0001000001100010111101011100001001100101101000";
      when  905 => r := "0001000000111100011100011100001011101101110010";
      when  906 => r := "0001000000010101111111111100001101110101110110";
      when  907 => r := "0000111111101111100110111100001111111101110111";
      when  908 => r := "0000111111001001010010011100010010000101110010";
      when  909 => r := "0000111110100011000001011100010100001101101010";
      when  910 => r := "0000111101111100110100111100010110010101011011";
      when  911 => r := "0000111101010110101100011100011000011101001000";
      when  912 => r := "0000111100110000100111011100011010100100110010";
      when  913 => r := "0000111100001010100110111100011100101100010101";
      when  914 => r := "0000111011100100101010011100011110110011110011";
      when  915 => r := "0000111010111110110001111100100000111011001101";
      when  916 => r := "0000111010011000111100111100100011000010100100";
      when  917 => r := "0000111001110011001100011100100101001001110100";
      when  918 => r := "0000111001001101011111011100100111010001000001";
      when  919 => r := "0000111000100111110110111100101001011000000111";
      when  920 => r := "0000111000000010010001111100101011011111001010";
      when  921 => r := "0000110111011100110000111100101101100110001000";
      when  922 => r := "0000110110110111010011111100101111101101000001";
      when  923 => r := "0000110110010001111010011100110001110011110110";
      when  924 => r := "0000110101101100100101011100110011111010100101";
      when  925 => r := "0000110101000111010011111100110110000001010001";
      when  926 => r := "0000110100100010000110011100111000000111110111";
      when  927 => r := "0000110011111100111100011100111010001110011010";
      when  928 => r := "0000110011010111110110011100111100010100111000";
      when  929 => r := "0000110010110010110100011100111110011011010000";
      when  930 => r := "0000110010001101110110011101000000100001100011";
      when  931 => r := "0000110001101000111011111101000010100111110011";
      when  932 => r := "0000110001000100000101011101000100101101111101";
      when  933 => r := "0000110000011111010010011101000110110100000100";
      when  934 => r := "0000101111111010100011011101001000111010000110";
      when  935 => r := "0000101111010101111000011101001011000000000010";
      when  936 => r := "0000101110110001010000111101001101000101111010";
      when  937 => r := "0000101110001100101100111101001111001011101111";
      when  938 => r := "0000101101101000001100111101010001010001011110";
      when  939 => r := "0000101101000011110000011101010011010111001010";
      when  940 => r := "0000101100011111010111111101010101011100110000";
      when  941 => r := "0000101011111011000011011101010111100010010000";
      when  942 => r := "0000101011010110110001111101011001100111101111";
      when  943 => r := "0000101010110010100100011101011011101101000111";
      when  944 => r := "0000101010001110011010111101011101110010011010";
      when  945 => r := "0000101001101010010100111101011111110111101001";
      when  946 => r := "0000101001000110010010011101100001111100110101";
      when  947 => r := "0000101000100010010011011101100100000001111100";
      when  948 => r := "0000100111111110011000011101100110000110111101";
      when  949 => r := "0000100111011010100000111101101000001011111011";
      when  950 => r := "0000100110110110101100111101101010010000110100";
      when  951 => r := "0000100110010010111100011101101100010101101010";
      when  952 => r := "0000100101101111001111111101101110011010011001";
      when  953 => r := "0000100101001011100110111101110000011111000101";
      when  954 => r := "0000100100101000000001011101110010100011101100";
      when  955 => r := "0000100100000100011111011101110100101000001111";
      when  956 => r := "0000100011100001000000111101110110101100101110";
      when  957 => r := "0000100010111101100110011101111000110001000111";
      when  958 => r := "0000100010011010001110111101111010110101011101";
      when  959 => r := "0000100001110110111011011101111100111001101101";
      when  960 => r := "0000100001010011101011011101111110111101111001";
      when  961 => r := "0000100000110000011110011110000001000010000011";
      when  962 => r := "0000100000001101010101011110000011000110000110";
      when  963 => r := "0000011111101010001111111110000101001010000101";
      when  964 => r := "0000011111000111001101011110000111001110000010";
      when  965 => r := "0000011110100100001110111110001001010001111000";
      when  966 => r := "0000011110000001010011111110001011010101101001";
      when  967 => r := "0000011101011110011011111110001101011001011000";
      when  968 => r := "0000011100111011100111111110001111011101000001";
      when  969 => r := "0000011100011000110110111110010001100000100111";
      when  970 => r := "0000011011110110001001011110010011100100001000";
      when  971 => r := "0000011011010011011111011110010101100111100101";
      when  972 => r := "0000011010110000111000111110010111101010111101";
      when  973 => r := "0000011010001110010101111110011001101110010001";
      when  974 => r := "0000011001101011110110011110011011110001100000";
      when  975 => r := "0000011001001001011001111110011101110100101100";
      when  976 => r := "0000011000100111000000111110011111110111110011";
      when  977 => r := "0000011000000100101011011110100001111010110110";
      when  978 => r := "0000010111100010011001011110100011111101110011";
      when  979 => r := "0000010111000000001010011110100110000000101110";
      when  980 => r := "0000010110011101111110111110101000000011100100";
      when  981 => r := "0000010101111011110110111110101010000110010110";
      when  982 => r := "0000010101011001110001111110101100001001000100";
      when  983 => r := "0000010100110111110000111110101110001011101011";
      when  984 => r := "0000010100010101110010011110110000001110010001";
      when  985 => r := "0000010011110011110111111110110010010000110001";
      when  986 => r := "0000010011010010000000011110110100010011001101";
      when  987 => r := "0000010010110000001011111110110110010101100110";
      when  988 => r := "0000010010001110011010111110111000010111111010";
      when  989 => r := "0000010001101100101101011110111010011010001001";
      when  990 => r := "0000010001001011000010111110111100011100010101";
      when  991 => r := "0000010000101001011011111110111110011110011100";
      when  992 => r := "0000010000000111110111111111000000100000011111";
      when  993 => r := "0000001111100110010111011111000010100010011110";
      when  994 => r := "0000001111000100111001111111000100100100011001";
      when  995 => r := "0000001110100011011111011111000110100110010000";
      when  996 => r := "0000001110000010001000111111001000101000000001";
      when  997 => r := "0000001101100000110100111111001010101001110000";
      when  998 => r := "0000001100111111100100011111001100101011011010";
      when  999 => r := "0000001100011110010110111111001110101101000000";
      when 1000 => r := "0000001011111101001100111111010000101110100001";
      when 1001 => r := "0000001011011100000101111111010010101111111111";
      when 1002 => r := "0000001010111011000001111111010100110001011001";
      when 1003 => r := "0000001010011010000001011111010110110010101110";
      when 1004 => r := "0000001001111001000011111111011000110011111111";
      when 1005 => r := "0000001001011000001001011111011010110101001101";
      when 1006 => r := "0000001000110111010010011111011100110110010101";
      when 1007 => r := "0000001000010110011110011111011110110111011001";
      when 1008 => r := "0000000111110101101101011111100000111000011010";
      when 1009 => r := "0000000111010100111111011111100010111001011000";
      when 1010 => r := "0000000110110100010100111111100100111010001111";
      when 1011 => r := "0000000110010011101100111111100110111011000101";
      when 1012 => r := "0000000101110011001000011111101000111011110101";
      when 1013 => r := "0000000101010010100110111111101010111100100010";
      when 1014 => r := "0000000100110010001000111111101100111101001001";
      when 1015 => r := "0000000100010001101101011111101110111101101110";
      when 1016 => r := "0000000011110001010101011111110000111110001101";
      when 1017 => r := "0000000011010000111111111111110010111110101011";
      when 1018 => r := "0000000010110000101101111111110100111111000010";
      when 1019 => r := "0000000010010000011110111111110110111111010110";
      when 1020 => r := "0000000001110000010010111111111000111111100110";
      when 1021 => r := "0000000001010000001001111111111010111111110010";
      when 1022 => r := "0000000000110000000011111111111100111111111010";
      when 1023 => r := "0000000000010000000000111111111110111111111110";
      when others => r := (others => '0');
    end case;
    return r;
  end table;

  constant m_Nan : std_logic_vector (31 downto 0) := x"fff00000";

  signal ret : std_logic_vector (31 downto 0) := (others => '0');
  signal sign : std_logic := '0';
  signal expr_t : std_logic_vector (8 downto 0) := (others => '0');
  signal expr : std_logic_vector (7 downto 0) := (others => '0');
  signal key : std_logic_vector (9 downto 0) := (others => '0');
  signal raw_ret : std_logic_vector (45 downto 0) := (others => '0');
  signal h_a : std_logic_vector (12 downto 0) := (others => '0');
  signal h_b : std_logic_vector (12 downto 0) := (others => '0');
  signal l_a : std_logic_vector (10 downto 0) := (others => '0');
  signal l_b : std_logic_vector (10 downto 0) := (others => '0');
  signal HH : std_logic_vector (25 downto 0) := (others => '0');
  signal HL : std_logic_vector (23 downto 0) := (others => '0');
  signal LH : std_logic_vector (23 downto 0) := (others => '0');
  signal mul0 : std_logic_vector (25 downto 0) := (others => '0');
  signal mul : std_logic_vector (22 downto 0) := (others => '0');
  signal x_expr : std_logic_vector (7 downto 0) := (others => '0');
  signal m_a : std_logic_vector (24 downto 0) := (others => '0');
  signal m_b : std_logic_vector (24 downto 0) := (others => '0');
  signal sum : std_logic_vector (25 downto 0) := (others => '0');

begin  -- architecture rtl

  sign <= A (31);
  key <= (not A (23)) &  A(22 downto 14);
  expr_t <= "001111111" + A (30 downto 23);
  expr <= expr_t(8 downto 1);

  raw_ret <= table (key);

  h_a <= '1' & raw_ret (45 downto 34);
  h_b <= '1' & A (22 downto 11);
  l_a <= raw_ret (33 downto 23);
  l_b <= A (10 downto 0);

  HH <= h_a * h_b;
  HL <= h_a * l_b;
  LH <= l_a * h_b;

  mul0 <= "00000000000000000000000000" + HH + LH (23 downto 11) + HL (23 downto 11) + "10";

  with mul0 (25) select
    mul <=
    mul0 (24 downto 2) when '1',
    mul0 (23 downto 1) when others;

  x_expr <= x"81" when mul0 (25) = '1' and A (23) = '0' else
            x"80" when mul0 (25) = '1' or A (23) = '0' else
            x"7f";
          

  with x_expr select
    m_a <=
    "01" & mul (22 downto 0)      when x"7f",
    '1' & mul (22 downto 0) & '0' when others;

  with x_expr select
    m_b <=
    "01" & raw_ret (22 downto 0) when x"81",
    '1' & raw_ret (22 downto 0) & '0' when others;


  sum <= "00000000000000000000000000" + m_a + m_b;

  ret <= A when sign = '1' and A (30 downto 23) = x"00" else
         m_Nan when sign = '1' else
         x"00000000" when A (30 downto 23) = x"00" else
         A when A (30 downto 23) = x"ff" else
         sign & expr & sum (24 downto 2) when m_b (24) = '1' else
         sign & expr & sum (23 downto 1);  

  -- purpose: set ret -> Q
  -- type   : combinational
  -- inputs : CLK
  -- outputs: Q
  set_loop: process (CLK) is
  begin  -- process set_loop
    if rising_edge (CLK) then
      Q <= ret;
    end if;
  end process set_loop;


end architecture rtl;
