library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity fmul_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity fmul_tb;

architecture testbench of fmul_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "01000011000000000000000000000000",
    1 => "01000001101000000000000000000000",
    2 => "00111111000000000000000000000000",
    3 => "00111110001100101011100000000000",
    4 => "00111101001010101010011111011111",
    5 => "00111100011011100100011011000010",
    6 => "00111011101001100101100001110101",
    7 => "00111010111010000100001000100001",
    8 => "00111010101100111001000110010010",
    9 => "00111001111110101011100010001111",
    10 => "00111001001011110000100010000111",
    11 => "00111000011101000110001101110111",
    12 => "00110111101010101001110011001111",
    13 => "00110110111011100011011101010000",
    14 => "00111110001010101010101011000001",
    15 => "00111101011011100100101011001001",
    16 => "00111100101001100101101101000100",
    17 => "00111100000010001000011100100011",
    18 => "00111011001111101010000000101101",
    19 => "00111010100001010001010001100010",
    20 => "00111001101110011100111110100100",
    21 => "00111001000000011011011111101100",
    22 => "00111001010011011000010101011001",
    23 => "00111000100011110111101001101111",
    24 => "00110111110010000101010010000001",
    25 => "00110111000010111101101010111101",
    26 => "00110110010000110100010100111000",
    27 => "00110101100010000101001001111010",
    28 => "00110100101111100101011010100111",
    29 => "01000001111100000000000000000000",
    30 => "00111111000000000000000000000000",
    31 => "00111110100001100000101000000000",
    32 => "00111101001010101010011111011111",
    33 => "00111100101100101011010100010001",
    34 => "00111100001110110010001110000011",
    35 => "00111011110000111111011111001011",
    36 => "00111010101100111001000110010010",
    37 => "00111010001111000000101001101011",
    38 => "00111001110001001110100110011000",
    39 => "00111001010011100011001111101100",
    40 => "00111000110101111110111001110110",
    41 => "00111000011000100001111010000000",
    42 => "00111110001010101010101011000001",
    43 => "00111101101100101011100000010110",
    44 => "00111101001110110010011010101100",
    45 => "00111100000010001000011100100011",
    46 => "00111011100011101111100000100010",
    47 => "00111011000101011011011011101110",
    48 => "00111010100111001100011100110011",
    49 => "00111010001001000010110011001000",
    50 => "00111001010011011000010101011001",
    51 => "00111000110101110011011110100110",
    52 => "00111000011000010101111100010001",
    53 => "00110111111011000000000100100000",
    54 => "00110111011101110010001110011100",
    55 => "00110111000000010110011001001010",
    56 => "00110110100001111000000100110000",
    57 => "00111111011100001000111111010100",
    58 => "00111110111100001000111011100011",
    59 => "00111110101011110001110010001100",
    60 => "00111111011100001000111111010100",
    61 => "00111111010100000101010101101101",
    62 => "10111110101011110001110010001100",
    63 => "10111110101011110001110010001100",
    64 => "01000010010010000000000000000000",
    65 => "00111111000000000000000000000000",
    66 => "00111110101100101011100110110011",
    67 => "00111101001010101010011111011111",
    68 => "00111100111011100100100100000110",
    69 => "00111100101001100101101110011110",
    70 => "00111100011010000100100011000000",
    71 => "00111010101100111001000110010010",
    72 => "00111010011110101011101011110001",
    73 => "00111010001011110000101111011011",
    74 => "00111001111101000110101001101111",
    75 => "00111001101010101010001101001100",
    76 => "00111001011011100100001010100011",
    77 => "01000010010010000000000000000000",
    78 => "00111110001010101010101011000001",
    79 => "00111101111011100100110100001101",
    80 => "00111101101001100101111001101110",
    81 => "00111100000010001000011100100011",
    82 => "00111011101111101010000111111110",
    83 => "00111011100001010001011011101010",
    84 => "00111011001110011101010011110010",
    85 => "00111011000000011011110011011100",
    86 => "00111001010011011000010101011001",
    87 => "00111001000011110111101111001100",
    88 => "00111000110010000101100001010000",
    89 => "00111000100010111101111010111011",
    90 => "00111000010000110100110010100111",
    91 => "00111000000010000101100011110110",
    92 => "00110111101111100110000110000100",
    93 => "00111111000000000000000000000000",
    94 => "00111110101100101011100110110011",
    95 => "00111101001010101010011111011111",
    96 => "00111100111011100100100100000110",
    97 => "00111100101001100101101110011110",
    98 => "00111100011010000100100011000000",
    99 => "00111010101100111001000110010010",
    100 => "00111010011110101011101011110001",
    101 => "00111010001011110000101111011011",
    102 => "00111001111101000110101001101111",
    103 => "00111001101010101010001101001100",
    104 => "00111001011011100100001010100011",
    105 => "00111111001001001000111001110000",
    106 => "00111110001010101010101011000001",
    107 => "00111101111011100100110100001101",
    108 => "00111101101001100101111001101110",
    109 => "00111100000010001000011100100011",
    110 => "00111011101111101010000111111110",
    111 => "00111011100001010001011011101010",
    112 => "00111011001110011101010011110010",
    113 => "00111011000000011011110011011100",
    114 => "00111001010011011000010101011001",
    115 => "00111001000011110111101111001100",
    116 => "00111000110010000101100001010000",
    117 => "00111000100010111101111010111011",
    118 => "00111000010000110100110010100111",
    119 => "00111000000010000101100011110110",
    120 => "00110111101111100110000110000100",
    121 => "00111111001001001000111001110000",
    122 => "01000001110010000000000000000000",
    123 => "00111111100000000000000000000000",
    124 => "01000010001000000000000000000000",
    125 => "00111111100000000000000000000000",
    126 => "01000010100011000000000000000000",
    127 => "00111111100000000000000000000000",
    128 => "01000001111100000000000000000000",
    129 => "00111111100000000000000000000000",
    130 => "01000001111100000000000000000000",
    131 => "00111111100000000000000000000000",
    132 => "00000000000000000000000000000000",
    133 => "10111111110000000000000000000000",
    134 => "10111111100000000000000000000000",
    135 => "00000000000000000000000000000000",
    136 => "10111111110000000000000000000000",
    137 => "10111111100000000000000000000000",
    138 => "01000010001000000000000000000000",
    139 => "00111111100000000000000000000000",
    140 => "01000001111000000000000000000000",
    141 => "00111111100000000000000000000000",
    142 => "01000001111000000000000000000000",
    143 => "00111111100000000000000000000000",
    144 => "01000001011100000000000000000000",
    145 => "00111111100000000000000000000000",
    146 => "01000001011100000000000000000000",
    147 => "00111111100000000000000000000000",
    148 => "01000001011100000000000000000000",
    149 => "00111111100000000000000000000000",
    150 => "01000001110010000000000000000000",
    151 => "00111111100000000000000000000000",
    152 => "01000001110010000000000000000000",
    153 => "00111111100000000000000000000000",
    154 => "01000001111100000000000000000000",
    155 => "00111111100000000000000000000000",
    156 => "01000010001101000000000000000000",
    157 => "00111111100000000000000000000000",
    158 => "01000010100101100000000000000000",
    159 => "00111111100000000000000000000000",
    160 => "01000001110010000000000000000000",
    161 => "00111111100000000000000000000000",
    162 => "01000001001000000000000000000000",
    163 => "00111111100000000000000000000000",
    164 => "01000001001000000000000000000000",
    165 => "00111111100000000000000000000000",
    166 => "01000001110010000000000000000000",
    167 => "00111111100000000000000000000000",
    168 => "01000001101000000000000000000000",
    169 => "00111111100000000000000000000000",
    170 => "01000001101000000000000000000000",
    171 => "00111111100000000000000000000000",
    172 => "01000001101000000000000000000000",
    173 => "00111111100000000000000000000000",
    174 => "01000001101000000000000000000000",
    175 => "00111111100000000000000000000000",
    176 => "01000001101000000000000000000000",
    177 => "00111111100000000000000000000000",
    178 => "00000000000000000000000000000000",
    179 => "10111111100000000000000000000000",
    180 => "00000000000000000000000000000000",
    181 => "10111111100000000000000000000000",
    182 => "01000001000100000000000000000000",
    183 => "00000000000000000000000000000000",
    184 => "00111100111100110000100000110101",
    185 => "10111101001110100000110100100110",
    186 => "10111110001001010000000010100000",
    187 => "00111110110101100101110110110100",
    188 => "00111111101001111000110101110011",
    189 => "00111110001010101010101011000001",
    190 => "10111100101100101011100100011010",
    191 => "00111011001110110010100011001101",
    192 => "00111100000010001000011100100011",
    193 => "10111010100011101111100011110010",
    194 => "00111001000101011011100010100010",
    195 => "10110111100111001100100111011111",
    196 => "00110110001001000011000010000011",
    197 => "00111001010011011000010101011001",
    198 => "10110111110101110011100011011111",
    199 => "00110110011000010110000110100001",
    200 => "10110100111011000000010100100110",
    201 => "00110011011101110010100100111010",
    202 => "10110010000000010110100111110111",
    203 => "00110000100001111000010111001111",
    204 => "00111111000000000000000000000000",
    205 => "10111101100001100000101011000011",
    206 => "00111101001010101010011111011111",
    207 => "10111011101100101011011000010101",
    208 => "00111010001110110010010110100011",
    209 => "10111000110000111111101100100001",
    210 => "00111010101100111001000110010010",
    211 => "10111001001111000000101101111100",
    212 => "00110111110001001110101111010100",
    213 => "10110110010011100011011101101111",
    214 => "00110100110101111111001101011101",
    215 => "10110011011000100010010011101100",
    216 => "00111110000001011010100011011000",
    217 => "10111110000001101101000000011011",
    218 => "10111101001010101000011010111111",
    219 => "00111100111100110000100000110101",
    220 => "10111101001111010101011011000010",
    221 => "10111110001001100101001000100100",
    222 => "00111110110101101000100000000010",
    223 => "00111111101001100011101101110000",
    224 => "00111111000000000000000000000000",
    225 => "00111110010011011100111111001001",
    226 => "00111101001010101010011111011111",
    227 => "00111100100010010011001011110000",
    228 => "00111011110111001001101001001011",
    229 => "00111011001100010101101010011011",
    230 => "00111010101100111001000110010010",
    231 => "00111010000100000101110101010001",
    232 => "00111001011010000001111111001100",
    233 => "00111000101110101001110111011101",
    234 => "00111000000101100000011111100001",
    235 => "00110111011100010011110000101001",
    236 => "00111110001010101010101011000001",
    237 => "00111101100010010011010101000010",
    238 => "00111100110111001001111000000110",
    239 => "00111100000010001000011100100011",
    240 => "00111011010110111000011000001110",
    241 => "00111010101100000111110010000110",
    242 => "00111010000011011110001011110110",
    243 => "00111001011001000010001111010001",
    244 => "00111001010011011000010101011001",
    245 => "00111000101001010011101010010111",
    246 => "00111000000001001101011000000110",
    247 => "00110111010101011001011001100111",
    248 => "00110110101010111011011011001100",
    249 => "00110110000010100000110011000000",
    250 => "00110101010111011111100010000100",
    251 => "00111111011010111001100000011100",
    252 => "01000000000101101000101101010010",
    253 => "00111111010000000001000101110111",
    254 => "00111100111100110000100000110101",
    255 => "10111101110100101000100100000100",
    256 => "10111110000100110011010100101010",
    257 => "00111111010000000110110110010110",
    258 => "00111111011010001000000110101110",
    259 => "00111110001010101010101011000001",
    260 => "10111100011110000000000111101011",
    261 => "00111010101101000011001010110010",
    262 => "00111100000010001000011100100011",
    263 => "10111010010001100110010111001110",
    264 => "00111000100100000010011100000010",
    265 => "10110110110100010111101000110010",
    266 => "00110101000110000011001111100010",
    267 => "00111001010011011000010101011001",
    268 => "10110111100101010101001111110111",
    269 => "00110101110110001111111110010100",
    270 => "10110100000111011010101011010101",
    271 => "00110010011001010001110111100110",
    272 => "10110000101001100111100011101101",
    273 => "00101110111100011110100101111000",
    274 => "00111111000000000000000000000000",
    275 => "10111101001110100000000101011001",
    276 => "00111101001010101010011111011111",
    277 => "10111011011101111111110110111011",
    278 => "00111001101101000010111110100111",
    279 => "10111000000000101110101110010001",
    280 => "00111010101100111001000110010010",
    281 => "10111001000000100111100010110101",
    282 => "00110111001111011001100011000110",
    283 => "10110101100010011100000111111111",
    284 => "00110011110010000010111101011001",
    285 => "10110010000100010111001101110011",
    286 => "00111101101110011011111111101000",
    287 => "10111101101110101000010010110101",
    288 => "10111101100101111101110001011011",
    289 => "00111100111100110000100000110101",
    290 => "10111101010001000011001011110000",
    291 => "10111110001010001110110111000100",
    292 => "00111110110101110011011000100010",
    293 => "00111111101000111011101001011000",
    294 => "00111111000000000000000000000000",
    295 => "00111110010101101101001110111001",
    296 => "00111101001010101010011111011111",
    297 => "00111100100011110011010101110111",
    298 => "00111011111100000101101001000011",
    299 => "00111011010010011011001000111011",
    300 => "00111010101100111001000110010010",
    301 => "00111010000101101011000000110010",
    302 => "00111001011111001110011111010011",
    303 => "00111000110101000011101011110011",
    304 => "00111000001100100001100011001100",
    305 => "00110111100101010111010000000101",
    306 => "00111110001010101010101011000001",
    307 => "00111101100011110011011111100011",
    308 => "00111100111100000101111001010011",
    309 => "00111100000010001000011100100011",
    310 => "00111011011001010010001111000010",
    311 => "00111010110000000100100101100101",
    312 => "00111010001000010101110001100001",
    313 => "00111001100001110110100010101100",
    314 => "00111001010011011000010101011001",
    315 => "00111000101011000111011101110001",
    316 => "00111000000100001011101001111011",
    317 => "00110111011100101110011100101001",
    318 => "00110110110010111101011000011111",
    319 => "00110110001010110000110110010010",
    320 => "00110101100011111000101011001111",
    321 => "00111111011010011100101101001110",
    322 => "01000000000011110111100101011101",
    323 => "00111111001110100110011110001000",
    324 => "00111100111100110000100000110101",
    325 => "10111101110100001001111110000100",
    326 => "10111110000101010101000011110010",
    327 => "00111111001111101001101100011010",
    328 => "00111111011011000100010001011010",
    329 => "00111110001010101010101011000001",
    330 => "10111100011111000000010011000101",
    331 => "00111010101110100001001011110010",
    332 => "00111100000010001000011100100011",
    333 => "10111010010010011001101101000000",
    334 => "00111000100101001101101001011100",
    335 => "10110110110110111100111001111000",
    336 => "00110101001000100100101001101011",
    337 => "00111001010011011000010101011001",
    338 => "10110111100101111011111000111110",
    339 => "00110101111000000001001100001000",
    340 => "10110100001001010111000100011001",
    341 => "00110010011101000100110101111111",
    342 => "10110000101101000110000010001001",
    343 => "00101111000001010010110110111001",
    344 => "00111111000000000000000000000000",
    345 => "10111101001111010000001101111100",
    346 => "00111101001010101010011111011111",
    347 => "10111011011111000000000010000011",
    348 => "00111001101110100000111111001110",
    349 => "10111000000010010110000000110010",
    350 => "00111010101100111001000110010010",
    351 => "10111001000001001001010011101010",
    352 => "00110111010000111100011101111101",
    353 => "10110101100100001000110011110001",
    354 => "00110011110101010111010000001010",
    355 => "10110010000111011001100110010010",
    356 => "00111101101111001011111011010001",
    357 => "10111101101111011000110101010011",
    358 => "10111101100101100111100110011111",
    359 => "00111100111100110000100000110101",
    360 => "10111101010001000000010110010000",
    361 => "10111110001010001101110100100100",
    362 => "00111110110101110011000000110010",
    363 => "00111111101000111100100111011101",
    364 => "00111111000000000000000000000000",
    365 => "00111110010101101001101111011101",
    366 => "00111101001010101010011111011111",
    367 => "00111100100011110001000000111011",
    368 => "00111011111011111101110101010110",
    369 => "00111011010010010001010100001111",
    370 => "00111010101100111001000110010010",
    371 => "00111010000101101000100100000011",
    372 => "00111001011111000110010001011110",
    373 => "00111000110100111001010110010000",
    374 => "00111000001100010101111111010111",
    375 => "00110111100101001011001000011011",
    376 => "00111110001010101010101011000001",
    377 => "00111101100011110001001010100101",
    378 => "00111100111011111110000101100010",
    379 => "00111100000010001000011100100011",
    380 => "00111011011001001110100000101101",
    381 => "00111010101111111110010101110011",
    382 => "00111010001000001101111010100011",
    383 => "00111001100001101101110000001101",
    384 => "00111001010011011000010101011001",
    385 => "00111000101011000100101010011001",
    386 => "00111000000100000110111101000001",
    387 => "00110111011100100010100111100000",
    388 => "00110110110010110000001001110001",
    389 => "00110110001010100010111110100011",
    390 => "00110101100011101010101101101111",
    391 => "00111111011010011101011010101110",
    392 => "01000000000011111010001101111010",
    393 => "00111111001110101000011110100001",
    394 => "00111100111100110000100000110101",
    395 => "10111101110100001010101010011001",
    396 => "10111110000101010100010011100110",
    397 => "00111111001111101010010110110011",
    398 => "00111111011011000010111011110000",
    399 => "00111110001010101010101011000001",
    400 => "10111100011110111110110111101101",
    401 => "00111010101110011111000100111000",
    402 => "00111100000010001000011100100011",
    403 => "10111010010010011000100011111010",
    404 => "00111000100101001011111101100001",
    405 => "10110110110110111001001010111000",
    406 => "00110101001000100000111110011100",
    407 => "00111001010011011000010101011001",
    408 => "10110111100101111011000001111101",
    409 => "00110101110111111110101001101011",
    410 => "10110100001001010100010000100000",
    411 => "00110010011100111111010011110111",
    412 => "10110000101101000000111011011000",
    413 => "00101111000001001110010101011011",
    414 => "00111111000000000000000000000000",
    415 => "10111101001111001111001001011010",
    416 => "00111101001010101010011111011111",
    417 => "10111011011110111110100110101100",
    418 => "00111001101110011110111000010101",
    419 => "10111000000010010011101011011011",
    420 => "00111010101100111001000110010010",
    421 => "10111001000001001000100011100101",
    422 => "00110111010000111010010000000000",
    423 => "10110101100100000110010110100101",
    424 => "00110011110101010010011010101111",
    425 => "10110010000111010101001000110001",
    426 => "00111101101111001010110111000001",
    427 => "10111101101111010111110000001110",
    428 => "10111101100101101000000110110101",
    429 => "00111100111100110000100000110101",
    430 => "10111101010001000000011010011010",
    431 => "10111110001010001101110110000100",
    432 => "00111110110101110011000001011000",
    433 => "00111111101000111100100110000101",
    434 => "00111111000000000000000000000000",
    435 => "00111110010101101001110100011001",
    436 => "00111101001010101010011111011111",
    437 => "00111100100011110001000100001101",
    438 => "00111011111011111110000000010111",
    439 => "00111011010010010001100010000110",
    440 => "00111010101100111001000110010010",
    441 => "00111010000101101000100111100001",
    442 => "00111001011111000110011101000110",
    443 => "00111000110100111001100100110111",
    444 => "00111000001100010110001111101101",
    445 => "00110111100101001011011001100011",
    446 => "00111110001010101010101011000001",
    447 => "00111101100011110001001101111000",
    448 => "00111100111011111110010000100101",
    449 => "00111100000010001000011100100011",
    450 => "00111011011001001110100101111110",
    451 => "00111010101111111110011110101000",
    452 => "00111010001000001110000101101001",
    453 => "00111001100001101101111100100111",
    454 => "00111001010011011000010101011001",
    455 => "00111000101011000100101110010110",
    456 => "00111000000100000111000011101010",
    457 => "00110111011100100010111000001101",
    458 => "00110110110010110000011100011011",
    459 => "00110110001010100011010010000111",
    460 => "00110101100011101011000001011011",
    461 => "00111111011010011101011001101110",
    462 => "01000000000011111010001010001011",
    463 => "00111111001110101000011011101101",
    464 => "00111100111100110000100000110101",
    465 => "10111101110100001010101001011010",
    466 => "10111110000101010100010100101010",
    467 => "00111111001111101010010101111000",
    468 => "00111111011011000010111101101010",
    469 => "00111110001010101010101011000001",
    470 => "10111100011110111110111001110000",
    471 => "00111010101110011111000111111010",
    472 => "00111100000010001000011100100011",
    473 => "10111010010010011000100101100010",
    474 => "00111000100101001011111111111011",
    475 => "10110110110110111001010000001101",
    476 => "00110101001000100001000011101100",
    477 => "00111001010011011000010101011001",
    478 => "10110111100101111011000011001011",
    479 => "00110101110111111110101101010010",
    480 => "10110100001001010100010100100000",
    481 => "00110010011100111111011011101111",
    482 => "10110000101101000001000010101001",
    483 => "00101111000001001110011011110111",
    484 => "00111111000000000000000000000000",
    485 => "10111101001111001111001010111100",
    486 => "00111101001010101010011111011111",
    487 => "10111011011110111110101000101110",
    488 => "00111001101110011110111011010101",
    489 => "10111000000010010011101110110000",
    490 => "00111010101100111001000110010010",
    491 => "10111001000001001000100100101010",
    492 => "00110111010000111010010011001011",
    493 => "10110101100100000110011010000110",
    494 => "00110011110101010010100001101010",
    495 => "10110010000111010101001111001010",
    496 => "00111101101111001010111000100011",
    497 => "10111101101111010111110001110000",
    498 => "10111101100101101000000110001000",
    499 => "00111100111100110000100000110101",
    500 => "10111101010001000000011010010010",
    501 => "10111110001010001101110110000010",
    502 => "00111110110101110011000001010110",
    503 => "00111111101000111100100110000110",
    504 => "00111111000000000000000000000000",
    505 => "00111110010101101001110100010101",
    506 => "00111101001010101010011111011111",
    507 => "00111100100011110001000100001010",
    508 => "00111011111011111110000000001110",
    509 => "00111011010010010001100001111011",
    510 => "00111010101100111001000110010010",
    511 => "00111010000101101000100111011110",
    512 => "00111001011111000110011100111100",
    513 => "00111000110100111001100100101011",
    514 => "00111000001100010110001111011111",
    515 => "00110111100101001011011001010100",
    516 => "00111110001010101010101011000001",
    517 => "00111101100011110001001101110101",
    518 => "00111100111011111110010000011100",
    519 => "00111100000010001000011100100011",
    520 => "00111011011001001110100101111001",
    521 => "00111010101111111110011110100000",
    522 => "00111010001000001110000101100000",
    523 => "00111001100001101101111100011101",
    524 => "00111001010011011000010101011001",
    525 => "00111000101011000100101110010011",
    526 => "00111000000100000111000011100101",
    527 => "00110111011100100010111000000000",
    528 => "00110110110010110000011100001101",
    529 => "00110110001010100011010001111000",
    530 => "00110101100011101011000001001011",
    531 => "00111111011010011101011001101110",
    532 => "01000000000011111010001010001101",
    533 => "10111101100101101000000110001000",
    534 => "00111111001110101000011011101101",
    535 => "10111101100101101000000110001000",
    536 => "00111111001110101000011011101101",
    537 => "00000000000000000000000000000000",
    538 => "00111100111100110000100000110101",
    539 => "10111101001110100000110100100110",
    540 => "10111110001001010000000010100000",
    541 => "00111110110101100101110110110100",
    542 => "00111111101001111000110101110011",
    543 => "00111111000000000000000000000000",
    544 => "00111110010010010000111011111001",
    545 => "00111101001010101010011111011111",
    546 => "00111100100001100000011111001000",
    547 => "00111011110100101000011111100101",
    548 => "00111011001001010101100100000010",
    549 => "00111010101100111001000110010010",
    550 => "00111010000011010000011111001011",
    551 => "00111001010111011000011010111011",
    552 => "00111000101011011111101110111101",
    553 => "00111000000010001010010011010100",
    554 => "00110111010101101010001011010000",
    555 => "00111110001010101010101011000001",
    556 => "00111101100001100000101000001100",
    557 => "00111100110100101000101101110100",
    558 => "00111100000010001000011100100011",
    559 => "00111011010101100111010000101100",
    560 => "00111010101010000110110111000000",
    561 => "00111010000001000100100000000101",
    562 => "00111001010011111100100010010000",
    563 => "00111001010011011000010101011001",
    564 => "00111000101000010110100110110111",
    565 => "00110111111111011000101011100010",
    566 => "00110111010001110010000011011111",
    567 => "00110110100111000110010001110100",
    568 => "00110101111101011010100000001000",
    569 => "00110101010000001110111101001011",
    570 => "00111111011011001000001110001010",
    571 => "01000000000110101000001100111110",
    572 => "00111111010000110111000111011101",
    573 => "00111100111100110000100000110101",
    574 => "10111101110100111010001001011110",
    575 => "10111110000100011111011111110010",
    576 => "00111111010000010111011111111001",
    577 => "00111111011001100100100011111000",
    578 => "00111111000000000000000000000000",
    579 => "00111110110000101101111000000100",
    580 => "00111101001010101010011111011111",
    581 => "00111101000000011110011100110110",
    582 => "00111100110001011100001110111110",
    583 => "00111100100101101000100111011000",
    584 => "00111010101100111001000110010010",
    585 => "00111010100010001011000000001011",
    586 => "00111010010100000001011111100101",
    587 => "00111010000111100110011010010010",
    588 => "00111001111100010010011000110011",
    589 => "00111001101101111001000000010100",
    590 => "00111110001010101010101011000001",
    591 => "00111110000000011110100101101000",
    592 => "00111101110001011100011100010101",
    593 => "00111100000010001000011100100011",
    594 => "00111011110011111101100110011111",
    595 => "00111011100111100011011100101011",
    596 => "00111011011100001101111000001000",
    597 => "00111011001101110101100100100101",
    598 => "00111001010011011000010101011001",
    599 => "00111001000111000111000101001001",
    600 => "00111000111011100010101100001011",
    601 => "00111000101101010100101100101010",
    602 => "00111000100010100000000000101111",
    603 => "00111000010100100001011110100011",
    604 => "00111000000111111110110000011100",
    605 => "00111111001110010101100010100010",
    606 => "00111111100001100101100110000001",
    607 => "00111111010111100000101010011001",
    608 => "00111100111100110000100000110101",
    609 => "10111101110110110101100011001100",
    610 => "10111110000010001011011010010111",
    611 => "00111111010010001001101101110110",
    612 => "00111111010101010111010101101100",
    613 => "00111110001010101010101011000001",
    614 => "00111110000000000001001101010001",
    615 => "00111101110000000011100111011111",
    616 => "00111100000010001000011100100011",
    617 => "00111011110011001110100110000010",
    618 => "00111011100110011100011000111111",
    619 => "00111011011001101100110000010000",
    620 => "00111011001011010011001100010101",
    621 => "00111001010011011000010101011001",
    622 => "00111001000110100011101100110010",
    623 => "00111000111001110111101110010111",
    624 => "00111000101011011011011011001110",
    625 => "00111000100000100101110010110011",
    626 => "00111000010000111010100001110110",
    627 => "00111000000100101101010001101011",
    628 => "00111111000000000000000000000000",
    629 => "00111110110000000001110011100010",
    630 => "00111101001010101010011111011111",
    631 => "00111101000000000001000100100111",
    632 => "00111100110000000011011010100000",
    633 => "00111100100100000011111010100111",
    634 => "00111010101100111001000110010010",
    635 => "00111010100001101100000101101111",
    636 => "00111010010010100100000010001110",
    637 => "00111010000101111100011100111011",
    638 => "00111001111000111100110100010111",
    639 => "00111001101010101111001110000100",
    640 => "00111111001011101001010011111111",
    641 => "00111111011011101011001100010011",
    642 => "00111111010111000101110111101110",
    643 => "00111100111100110000100000110101",
    644 => "10111101110110101110011111110010",
    645 => "10111110000010010100010011000010",
    646 => "00111111010010000011010100111001",
    647 => "00111111010101100111101010000110",
    648 => "00111110001010101010101011000001",
    649 => "00111110000000001010111111111011",
    650 => "00111101110000100001000101000011",
    651 => "00111100000010001000011100100011",
    652 => "00111011110011011110010000101001",
    653 => "00111011100110110011111101011000",
    654 => "00111011011010100001111100010000",
    655 => "00111011001100001000100010011110",
    656 => "00111001010011011000010101011001",
    657 => "00111001000110101111011111011010",
    658 => "00111000111010011011001100111111",
    659 => "00111000101100000011011101010011",
    660 => "00111000100001001101111100100001",
    661 => "00111000010010000110000010011100",
    662 => "00111000000101110001011011111111",
    663 => "00111111000000000000000000000000",
    664 => "00111110110000010000011111100001",
    665 => "00111101001010101010011111011111",
    666 => "00111101000000001010110111001111",
    667 => "00111100110000100000110111111101",
    668 => "00111100100100100101001010000011",
    669 => "00111010101100111001000110010010",
    670 => "00111010100001110110011001000101",
    671 => "00111010010011000011000010001001",
    672 => "00111010000110011111011011011111",
    673 => "00111001111010000010111110110101",
    674 => "00111001101011110001001100011011",
    675 => "00111111001011110100000010010100",
    676 => "00111111011100000110101111010110",
    677 => "00111111010111000111101011001000",
    678 => "00111100111100110000100000110101",
    679 => "10111101110110101110111110010110",
    680 => "10111110000010010011101100101010",
    681 => "00111111010010000011110000100110",
    682 => "00111111010101100110100011101010",
    683 => "00111110001010101010101011000001",
    684 => "00111110000000001010010101101001",
    685 => "00111101110000011111000101100011",
    686 => "00111100000010001000011100100011",
    687 => "00111011110011011101001101000000",
    688 => "00111011100110110010010111011001",
    689 => "00111011011010011110010101100101",
    690 => "00111011001100000100111010100110",
    691 => "00111001010011011000010101011001",
    692 => "00111001000110101110101100100000",
    693 => "00111000111010011000110011011110",
    694 => "00111000101100000000101111101011",
    695 => "00111000100001001011001101111111",
    696 => "00111000010010000000111001100000",
    697 => "00111000000101101100110010011010",
    698 => "00111111000000000000000000000000",
    699 => "00111110110000001111100000000110",
    700 => "00111101001010101010011111011111",
    701 => "00111101000000001010001100111101",
    702 => "00111100110000011110111000011101",
    703 => "00111100100100100010111001111000",
    704 => "00111010101100111001000110010010",
    705 => "00111010100001110101101100100110",
    706 => "00111010010011000000111011111111",
    707 => "00111010000110011101000011110010",
    708 => "00111001111001111110001101110110",
    709 => "00111001101011101100101101000001",
    710 => "00111111001011110011010100000110",
    711 => "00111111011100000100111000001000",
    712 => "00111111010111000111100011011111",
    713 => "00111100111100110000100000110101",
    714 => "10111101110110101110111100010100",
    715 => "10111110000010010011101111001100",
    716 => "00111111010010000011101110110001",
    717 => "00111111010101100110101000010100",
    718 => "00111110001010101010101011000001",
    719 => "00111110000000001010011000011101",
    720 => "00111101110000011111001110000010",
    721 => "00111100000010001000011100100011",
    722 => "00111011110011011101010001100000",
    723 => "00111011100110110010011110001011",
    724 => "00111011011010011110100100111011",
    725 => "00111011001100000101001010000001",
    726 => "00111001010011011000010101011001",
    727 => "00111001000110101110101111111001",
    728 => "00111000111010011000111101101100",
    729 => "00111000101100000000111011001111",
    730 => "00111000100001001011011001100111",
    731 => "00111000010010000001001111011001",
    732 => "00111000000101101101000110001101",
    733 => "00111111000000000000000000000000",
    734 => "00111110110000001111100100010100",
    735 => "00111101001010101010011111011111",
    736 => "00111101000000001010001111110001",
    737 => "00111100110000011111000000111100",
    738 => "00111100100100100011000011011110",
    739 => "00111010101100111001000110010010",
    740 => "00111010100001110101101111100011",
    741 => "00111010010011000001000100111010",
    742 => "00111010000110011101001101110111",
    743 => "00111001111001111110100010000111",
    744 => "00111001101011101101000000001000",
    745 => "00111111001011110011010111001010",
    746 => "00111111011100000101000000000010",
    747 => "00111111010111000111100100000001",
    748 => "00111100111100110000100000110101",
    749 => "10111101110110101110111100011101",
    750 => "10111110000010010011101111000010",
    751 => "00111111010010000011101110111001",
    752 => "00111111010101100110101000000000",
    753 => "00111110001010101010101011000001",
    754 => "00111110000000001010011000010001",
    755 => "00111101110000011111001101011101",
    756 => "00111100000010001000011100100011",
    757 => "00111011110011011101010001001100",
    758 => "00111011100110110010011101101100",
    759 => "00111011011010011110100011110101",
    760 => "00111011001100000101001000111011",
    761 => "00111001010011011000010101011001",
    762 => "00111001000110101110101111101001",
    763 => "00111000111010011000111100111101",
    764 => "00111000101100000000111010011010",
    765 => "00111000100001001011011000110010",
    766 => "00111000010010000001001101110110",
    767 => "00111000000101101101000100110011",
    768 => "00111111000000000000000000000000",
    769 => "00111110110000001111100100000001",
    770 => "00111101001010101010011111011111",
    771 => "00111101000000001010001111100100",
    772 => "00111100110000011111000000010101",
    773 => "00111100100100100011000010110010",
    774 => "00111010101100111001000110010010",
    775 => "00111010100001110101101111010110",
    776 => "00111010010011000001000100010010",
    777 => "00111010000110011101001101001010",
    778 => "00111001111001111110100000101100",
    779 => "00111001101011101100111110110010",
    780 => "00111111001011110011010110111100",
    781 => "00111111011100000100111111011111",
    782 => "00111111010111000111100011111110",
    783 => "00111100111100110000100000110101",
    784 => "10111101110110101110111100011100",
    785 => "10111110000010010011101111000011",
    786 => "00111111010010000011101110111000",
    787 => "00111111010101100110101000000010",
    788 => "00111110001010101010101011000001",
    789 => "00111110000000001010011000010011",
    790 => "00111101110000011111001101100011",
    791 => "00111100000010001000011100100011",
    792 => "00111011110011011101010001001111",
    793 => "00111011100110110010011101110001",
    794 => "00111011011010011110100100000000",
    795 => "00111011001100000101001001000110",
    796 => "00111001010011011000010101011001",
    797 => "00111001000110101110101111101100",
    798 => "00111000111010011000111101000101",
    799 => "00111000101100000000111010100011",
    800 => "00111000100001001011011000111010",
    801 => "00111000010010000001001110000101",
    802 => "00111000000101101101000101000001",
    803 => "00111111000000000000000000000000",
    804 => "00111110110000001111100100000100",
    805 => "00111101001010101010011111011111",
    806 => "00111101000000001010001111100110",
    807 => "00111100110000011111000000011011",
    808 => "00111100100100100011000010111001",
    809 => "00111010101100111001000110010010",
    810 => "00111010100001110101101111011000",
    811 => "00111010010011000001000100011000",
    812 => "00111010000110011101001101010001",
    813 => "00111001111001111110100000111010",
    814 => "00111001101011101100111110111111",
    815 => "00111111001011110011010110111111",
    816 => "00111111011100000100111111100110",
    817 => "00111111010111000111100100000001",
    818 => "00111100111100110000100000110101",
    819 => "10111101110110101110111100011101",
    820 => "10111110000010010011101111000010",
    821 => "00111111010010000011101110111001",
    822 => "00111111010101100110101000000000",
    823 => "00111110001010101010101011000001",
    824 => "00111110000000001010011000010001",
    825 => "00111101110000011111001101011101",
    826 => "00111100000010001000011100100011",
    827 => "00111011110011011101010001001100",
    828 => "00111011100110110010011101101100",
    829 => "00111011011010011110100011110101",
    830 => "00111011001100000101001000111011",
    831 => "00111001010011011000010101011001",
    832 => "00111001000110101110101111101001",
    833 => "00111000111010011000111100111101",
    834 => "00111000101100000000111010011010",
    835 => "00111000100001001011011000110010",
    836 => "00111000010010000001001101110110",
    837 => "00111000000101101101000100110011",
    838 => "00111111000000000000000000000000",
    839 => "00111110110000001111100100000001",
    840 => "00111101001010101010011111011111",
    841 => "00111101000000001010001111100100",
    842 => "00111100110000011111000000010101",
    843 => "00111100100100100011000010110010",
    844 => "00111010101100111001000110010010",
    845 => "00111010100001110101101111010110",
    846 => "00111010010011000001000100010010",
    847 => "00111010000110011101001101001010",
    848 => "00111001111001111110100000101100",
    849 => "00111001101011101100111110110010",
    850 => "00111111001011110011010110111100",
    851 => "00111111011100000100111111011111",
    852 => "00111111010111000111100011111110",
    853 => "00111100111100110000100000110101",
    854 => "10111101110110101110111100011100",
    855 => "10111110000010010011101111000011",
    856 => "00111111010010000011101110111000",
    857 => "00111111010101100110101000000010",
    858 => "00111110001010101010101011000001",
    859 => "00111110000000001010011000010011",
    860 => "00111101110000011111001101100011",
    861 => "00111100000010001000011100100011",
    862 => "00111011110011011101010001001111",
    863 => "00111011100110110010011101110001",
    864 => "00111011011010011110100100000000",
    865 => "00111011001100000101001001000110",
    866 => "00111001010011011000010101011001",
    867 => "00111001000110101110101111101100",
    868 => "00111000111010011000111101000101",
    869 => "00111000101100000000111010100011",
    870 => "00111000100001001011011000111010",
    871 => "00111000010010000001001110000101",
    872 => "00111000000101101101000101000001",
    873 => "00111111000000000000000000000000",
    874 => "00111110110000001111100100000100",
    875 => "00111101001010101010011111011111",
    876 => "00111101000000001010001111100110",
    877 => "00111100110000011111000000011011",
    878 => "00111100100100100011000010111001",
    879 => "00111010101100111001000110010010",
    880 => "00111010100001110101101111011000",
    881 => "00111010010011000001000100011000",
    882 => "00111010000110011101001101010001",
    883 => "00111001111001111110100000111010",
    884 => "00111001101011101100111110111111",
    885 => "00111111001011110011010110111111",
    886 => "00111111011100000100111111100110",
    887 => "00111111010111000111100011111110",
    888 => "00111111010111000111100100000001",
    889 => "00111111010111000111100011111110",
    890 => "00111111010111000111100100000001",
    891 => "01000000010000000000000000000000",
    892 => "00000000000000000000000000000000",
    893 => "00111100111100110000100000110101",
    894 => "10111101001110100000110100100110",
    895 => "10111110001001010000000010100000",
    896 => "00111110110101100101110110110100",
    897 => "00111111101001111000110101110011",
    898 => "00111110001010101010101011000001",
    899 => "10111101100001100000101011010011",
    900 => "00111100110100101000110111100101",
    901 => "00111100000010001000011100100011",
    902 => "10111011010101100111010101101010",
    903 => "00111010101010000110111110110100",
    904 => "10111010000001000100101001010010",
    905 => "00111001010011111100110101100010",
    906 => "00111001010011011000010101011001",
    907 => "10111000101000010110101010100110",
    908 => "00110111111111011000110111010001",
    909 => "10110111010001110010010001010011",
    910 => "00110110100111000110100000010010",
    911 => "10110101111101011010111100100011",
    912 => "00110101010000001111010111111110",
    913 => "00111111000000000000000000000000",
    914 => "10111110010010010001000000100011",
    915 => "00111101001010101010011111011111",
    916 => "10111100100001100000100010001111",
    917 => "00111011110100101000101001010110",
    918 => "10111011001001010101101111100010",
    919 => "00111010101100111001000110010010",
    920 => "10111010000011010000100010011100",
    921 => "00111001010111011000100101001100",
    922 => "10111000101011011111111011000011",
    923 => "00111000000010001010011111111110",
    924 => "10110111010101101010100100000110",
    925 => "00111110110000111110111101010110",
    926 => "10111110110101000001010000100000",
    927 => "10111110000001100010000101011011",
    928 => "00111100111100110000100000110101",
    929 => "10111101010101110100110101100010",
    930 => "10111110001011110010101110101110",
    931 => "00111110110110110101111100111000",
    932 => "00111111100111100100111011110111",
    933 => "00111111000000000000000000000000",
    934 => "00111110011010100101011001001101",
    935 => "00111101001010101010011111011111",
    936 => "00111100100111000011011011111001",
    937 => "00111100000011101111111011101000",
    938 => "00111011100000101110010100110100",
    939 => "00111010101100111001000110010010",
    940 => "00111010001001000101111110010111",
    941 => "00111001100101100111011011001001",
    942 => "00111001000010011011101101001100",
    943 => "00111000011111000010011101000010",
    944 => "00110111111001101101000011100010",
    945 => "00111110001010101010101011000001",
    946 => "00111101100111000011100110011100",
    947 => "00111101000011110000000101010010",
    948 => "00111100000010001000011100100011",
    949 => "00111011011110011111001100011000",
    950 => "00111010111001001100110001110110",
    951 => "00111010010100010111000000000100",
    952 => "00111001101111111011011011111101",
    953 => "00111001010011011000010101011001",
    954 => "00111000101111000010000100101011",
    955 => "00111000001011000011010110111100",
    956 => "00110111100111011010001100101011",
    957 => "00110111000100000100110001001001",
    958 => "00110110100001000001011001011111",
    959 => "00110101111100011101000111110011",
    960 => "00111111011001011010011011000011",
    961 => "01000000000000011110110111111101",
    962 => "00111111001100011110010000000101",
    963 => "00111100111100110000100000110101",
    964 => "10111101110011011001001110011100",
    965 => "10111110000110001000110100100110",
    966 => "00111111001110111010110010111100",
    967 => "00111111011100011111110000101100",
    968 => "00111110001010101010101011000001",
    969 => "10111101010000011001011010100010",
    970 => "00111100010110111001011010011000",
    971 => "00111100000010001000011100100011",
    972 => "10111011000110101101110100111110",
    973 => "00111010001011111010100111001010",
    974 => "10111001010001110100000101110010",
    975 => "00111000011000100000010001000010",
    976 => "00111001010011011000010101011001",
    977 => "10111000011010010001111110010010",
    978 => "00110111100001000011011101101001",
    979 => "10110110100101011111100101001000",
    980 => "00110101101010100001110110101111",
    981 => "10110100110000001111011010011101",
    982 => "00110011110110101110000100010101",
    983 => "00111111000000000000000000000000",
    984 => "10111110000100010011000011100111",
    985 => "00111101001010101010011111011111",
    986 => "10111100010000011001001101011101",
    987 => "00111011010110111001001011100011",
    988 => "10111010011110010001000001000111",
    989 => "00111010101100111001000110010010",
    990 => "10111001110010111010111110000001",
    991 => "00111000111001110000101010100000",
    992 => "10111000000000110000100100100110",
    993 => "00110111000101001010001001101100",
    994 => "10110110001010001001100011000111",
    995 => "00111110100011110100000010111101",
    996 => "10111110100101010011011001011010",
    997 => "10111110011000111101010110010001",
    998 => "00111100111100110000100000110101",
    999 => "10111101100000000000010111010001");

  constant b_lut : lut := (
    0 => "00111100000000000000000000000000",
    1 => "00111100100011101111100110011000",
    2 => "00111110101100101011011111111111",
    3 => "00111110101100101011011111111111",
    4 => "00111110101100101011011111111111",
    5 => "00111110101100101011011111111111",
    6 => "00111110101100101011011111111111",
    7 => "00111110101100101011011111111111",
    8 => "00111110101100101011011111111111",
    9 => "00111110101100101011011111111111",
    10 => "00111110101100101011011111111111",
    11 => "00111110101100101011011111111111",
    12 => "00111110101100101011011111111111",
    13 => "00111110101100101011011111111111",
    14 => "00111110101100101011011111111111",
    15 => "00111110101100101011011111111111",
    16 => "00111110101100101011011111111111",
    17 => "00111110101100101011011111111111",
    18 => "00111110101100101011011111111111",
    19 => "00111110101100101011011111111111",
    20 => "00111110101100101011011111111111",
    21 => "00111110101100101011011111111111",
    22 => "00111110101100101011011111111111",
    23 => "00111110101100101011011111111111",
    24 => "00111110101100101011011111111111",
    25 => "00111110101100101011011111111111",
    26 => "00111110101100101011011111111111",
    27 => "00111110101100101011011111111111",
    28 => "00111110101100101011011111111111",
    29 => "00111100100011101111100110011000",
    30 => "00111111000001100000100111111111",
    31 => "00111111000001100000100111111111",
    32 => "00111111000001100000100111111111",
    33 => "00111111000001100000100111111111",
    34 => "00111111000001100000100111111111",
    35 => "00111111000001100000100111111111",
    36 => "00111111000001100000100111111111",
    37 => "00111111000001100000100111111111",
    38 => "00111111000001100000100111111111",
    39 => "00111111000001100000100111111111",
    40 => "00111111000001100000100111111111",
    41 => "00111111000001100000100111111111",
    42 => "00111111000001100000100111111111",
    43 => "00111111000001100000100111111111",
    44 => "00111111000001100000100111111111",
    45 => "00111111000001100000100111111111",
    46 => "00111111000001100000100111111111",
    47 => "00111111000001100000100111111111",
    48 => "00111111000001100000100111111111",
    49 => "00111111000001100000100111111111",
    50 => "00111111000001100000100111111111",
    51 => "00111111000001100000100111111111",
    52 => "00111111000001100000100111111111",
    53 => "00111111000001100000100111111111",
    54 => "00111111000001100000100111111111",
    55 => "00111111000001100000100111111111",
    56 => "00111111000001100000100111111111",
    57 => "00111110111111111111111100000000",
    58 => "01000011010010000000000000000000",
    59 => "11000011010010000000000000000000",
    60 => "00111111010111011011010000100000",
    61 => "01000011010010000000000000000000",
    62 => "00111110111111111111111100000000",
    63 => "00111111010111011011010000100000",
    64 => "00111100100011101111100110011000",
    65 => "00111111001100101011100110110010",
    66 => "00111111001100101011100110110010",
    67 => "00111111001100101011100110110010",
    68 => "00111111001100101011100110110010",
    69 => "00111111001100101011100110110010",
    70 => "00111111001100101011100110110010",
    71 => "00111111001100101011100110110010",
    72 => "00111111001100101011100110110010",
    73 => "00111111001100101011100110110010",
    74 => "00111111001100101011100110110010",
    75 => "00111111001100101011100110110010",
    76 => "00111111001100101011100110110010",
    77 => "00111100100011101111100110011000",
    78 => "00111111001100101011100110110010",
    79 => "00111111001100101011100110110010",
    80 => "00111111001100101011100110110010",
    81 => "00111111001100101011100110110010",
    82 => "00111111001100101011100110110010",
    83 => "00111111001100101011100110110010",
    84 => "00111111001100101011100110110010",
    85 => "00111111001100101011100110110010",
    86 => "00111111001100101011100110110010",
    87 => "00111111001100101011100110110010",
    88 => "00111111001100101011100110110010",
    89 => "00111111001100101011100110110010",
    90 => "00111111001100101011100110110010",
    91 => "00111111001100101011100110110010",
    92 => "00111111001100101011100110110010",
    93 => "00111111001100101011100110110010",
    94 => "00111111001100101011100110110010",
    95 => "00111111001100101011100110110010",
    96 => "00111111001100101011100110110010",
    97 => "00111111001100101011100110110010",
    98 => "00111111001100101011100110110010",
    99 => "00111111001100101011100110110010",
    100 => "00111111001100101011100110110010",
    101 => "00111111001100101011100110110010",
    102 => "00111111001100101011100110110010",
    103 => "00111111001100101011100110110010",
    104 => "00111111001100101011100110110010",
    105 => "00111111010001000001101011100100",
    106 => "00111111001100101011100110110010",
    107 => "00111111001100101011100110110010",
    108 => "00111111001100101011100110110010",
    109 => "00111111001100101011100110110010",
    110 => "00111111001100101011100110110010",
    111 => "00111111001100101011100110110010",
    112 => "00111111001100101011100110110010",
    113 => "00111111001100101011100110110010",
    114 => "00111111001100101011100110110010",
    115 => "00111111001100101011100110110010",
    116 => "00111111001100101011100110110010",
    117 => "00111111001100101011100110110010",
    118 => "00111111001100101011100110110010",
    119 => "00111111001100101011100110110010",
    120 => "00111111001100101011100110110010",
    121 => "00111111001001001000111001110000",
    122 => "01000001110010000000000000000000",
    123 => "00111010110100011011011100010110",
    124 => "01000010001000000000000000000000",
    125 => "00111010001000111101011100001000",
    126 => "01000010100011000000000000000000",
    127 => "00111001010101011111111011000000",
    128 => "01000001111100000000000000000000",
    129 => "00111010100100011010001010110100",
    130 => "01000001111100000000000000000000",
    131 => "00111010100100011010001010110100",
    132 => "00000000000000000000000000000000",
    133 => "10111111110000000000000000000000",
    134 => "10111111100000000000000000000000",
    135 => "10111111000011100000000011010110",
    136 => "10111111000011100000000011010110",
    137 => "10111111000011100000000011010110",
    138 => "01000010001000000000000000000000",
    139 => "00111010001000111101011100001000",
    140 => "01000001111000000000000000000000",
    141 => "00111010101001110010111100000100",
    142 => "01000001111000000000000000000000",
    143 => "00111010101001110010111100000100",
    144 => "01000001011100000000000000000000",
    145 => "00111011100100011010001010110100",
    146 => "01000001011100000000000000000000",
    147 => "00111011100100011010001010110100",
    148 => "01000001011100000000000000000000",
    149 => "00111011100100011010001010110100",
    150 => "01000001110010000000000000000000",
    151 => "00111010110100011011011100010110",
    152 => "01000001110010000000000000000000",
    153 => "00111010110100011011011100010110",
    154 => "01000001111100000000000000000000",
    155 => "00111010100100011010001010110100",
    156 => "01000010001101000000000000000000",
    157 => "00111010000000010111010000101100",
    158 => "01000010100101100000000000000000",
    159 => "00111001001110100110100111011100",
    160 => "01000001110010000000000000000000",
    161 => "00111010110100011011011100010110",
    162 => "01000001001000000000000000000000",
    163 => "00111100001000111101011100001000",
    164 => "01000001001000000000000000000000",
    165 => "00111100001000111101011100001000",
    166 => "01000001110010000000000000000000",
    167 => "00111010110100011011011100010110",
    168 => "01000001101000000000000000000000",
    169 => "00111011001000111101011100001000",
    170 => "01000001101000000000000000000000",
    171 => "00111011001000111101011100001000",
    172 => "01000001101000000000000000000000",
    173 => "00111011001000111101011100001000",
    174 => "01000001101000000000000000000000",
    175 => "00111011001000111101011100001000",
    176 => "01000001101000000000000000000000",
    177 => "00111011001000111101011100001000",
    178 => "00000000000000000000000000000000",
    179 => "10111111100000000000000000000000",
    180 => "10111111100000000000000000000000",
    181 => "10111111100000000000000000000000",
    182 => "00111110010011001100110011001101",
    183 => "00000000000000000000000000000000",
    184 => "01000000010010100110001011000100",
    185 => "01000000010010100110001011000100",
    186 => "01000000010010100110001011000100",
    187 => "01000000010010100110001011000100",
    188 => "10111101110011001100110011001101",
    189 => "10111110000001100000101011000010",
    190 => "10111110000001100000101011000010",
    191 => "10111110000001100000101011000010",
    192 => "10111110000001100000101011000010",
    193 => "10111110000001100000101011000010",
    194 => "10111110000001100000101011000010",
    195 => "10111110000001100000101011000010",
    196 => "10111110000001100000101011000010",
    197 => "10111110000001100000101011000010",
    198 => "10111110000001100000101011000010",
    199 => "10111110000001100000101011000010",
    200 => "10111110000001100000101011000010",
    201 => "10111110000001100000101011000010",
    202 => "10111110000001100000101011000010",
    203 => "10111110000001100000101011000010",
    204 => "10111110000001100000101011000010",
    205 => "10111110000001100000101011000010",
    206 => "10111110000001100000101011000010",
    207 => "10111110000001100000101011000010",
    208 => "10111110000001100000101011000010",
    209 => "10111110000001100000101011000010",
    210 => "10111110000001100000101011000010",
    211 => "10111110000001100000101011000010",
    212 => "10111110000001100000101011000010",
    213 => "10111110000001100000101011000010",
    214 => "10111110000001100000101011000010",
    215 => "10111110000001100000101011000010",
    216 => "10111111100000010001101011000010",
    217 => "00111110101000011110100010011011",
    218 => "10111101001010101000011010111111",
    219 => "01000000010010001010011110000010",
    220 => "01000000010010001010011110000010",
    221 => "01000000010010001010011110000010",
    222 => "01000000010010001010011110000010",
    223 => "00111111011001100110011001101000",
    224 => "00111110110011011100111111001000",
    225 => "00111110110011011100111111001000",
    226 => "00111110110011011100111111001000",
    227 => "00111110110011011100111111001000",
    228 => "00111110110011011100111111001000",
    229 => "00111110110011011100111111001000",
    230 => "00111110110011011100111111001000",
    231 => "00111110110011011100111111001000",
    232 => "00111110110011011100111111001000",
    233 => "00111110110011011100111111001000",
    234 => "00111110110011011100111111001000",
    235 => "00111110110011011100111111001000",
    236 => "00111110110011011100111111001000",
    237 => "00111110110011011100111111001000",
    238 => "00111110110011011100111111001000",
    239 => "00111110110011011100111111001000",
    240 => "00111110110011011100111111001000",
    241 => "00111110110011011100111111001000",
    242 => "00111110110011011100111111001000",
    243 => "00111110110011011100111111001000",
    244 => "00111110110011011100111111001000",
    245 => "00111110110011011100111111001000",
    246 => "00111110110011011100111111001000",
    247 => "00111110110011011100111111001000",
    248 => "00111110110011011100111111001000",
    249 => "00111110110011011100111111001000",
    250 => "00111110110011011100111111001000",
    251 => "01000000001000111001010101100000",
    252 => "00111110101000110100111001000100",
    253 => "00111111010000000001000101110111",
    254 => "00111111100111010011011001010000",
    255 => "00111111100111010011011001010000",
    256 => "00111111100111010011011001010000",
    257 => "00111111100111010011011001010000",
    258 => "10111101110011001100110011001101",
    259 => "10111101101110100000000101011000",
    260 => "10111101101110100000000101011000",
    261 => "10111101101110100000000101011000",
    262 => "10111101101110100000000101011000",
    263 => "10111101101110100000000101011000",
    264 => "10111101101110100000000101011000",
    265 => "10111101101110100000000101011000",
    266 => "10111101101110100000000101011000",
    267 => "10111101101110100000000101011000",
    268 => "10111101101110100000000101011000",
    269 => "10111101101110100000000101011000",
    270 => "10111101101110100000000101011000",
    271 => "10111101101110100000000101011000",
    272 => "10111101101110100000000101011000",
    273 => "10111101101110100000000101011000",
    274 => "10111101101110100000000101011000",
    275 => "10111101101110100000000101011000",
    276 => "10111101101110100000000101011000",
    277 => "10111101101110100000000101011000",
    278 => "10111101101110100000000101011000",
    279 => "10111101101110100000000101011000",
    280 => "10111101101110100000000101011000",
    281 => "10111101101110100000000101011000",
    282 => "10111101101110100000000101011000",
    283 => "10111101101110100000000101011000",
    284 => "10111101101110100000000101011000",
    285 => "10111101101110100000000101011000",
    286 => "10111111100000001000011110011110",
    287 => "00111111010100000110111010001000",
    288 => "10111101100101111101110001011011",
    289 => "01000000010001010000101010010000",
    290 => "01000000010001010000101010010000",
    291 => "01000000010001010000101010010000",
    292 => "01000000010001010000101010010000",
    293 => "00111111011001100110011001101000",
    294 => "00111110110101101101001110111000",
    295 => "00111110110101101101001110111000",
    296 => "00111110110101101101001110111000",
    297 => "00111110110101101101001110111000",
    298 => "00111110110101101101001110111000",
    299 => "00111110110101101101001110111000",
    300 => "00111110110101101101001110111000",
    301 => "00111110110101101101001110111000",
    302 => "00111110110101101101001110111000",
    303 => "00111110110101101101001110111000",
    304 => "00111110110101101101001110111000",
    305 => "00111110110101101101001110111000",
    306 => "00111110110101101101001110111000",
    307 => "00111110110101101101001110111000",
    308 => "00111110110101101101001110111000",
    309 => "00111110110101101101001110111000",
    310 => "00111110110101101101001110111000",
    311 => "00111110110101101101001110111000",
    312 => "00111110110101101101001110111000",
    313 => "00111110110101101101001110111000",
    314 => "00111110110101101101001110111000",
    315 => "00111110110101101101001110111000",
    316 => "00111110110101101101001110111000",
    317 => "00111110110101101101001110111000",
    318 => "00111110110101101101001110111000",
    319 => "00111110110101101101001110111000",
    320 => "00111110110101101101001110111000",
    321 => "01000000000111010001100111101110",
    322 => "00111110101001100100110011011001",
    323 => "00111111001110100110011110001000",
    324 => "00111111101000010011110110001100",
    325 => "00111111101000010011110110001100",
    326 => "00111111101000010011110110001100",
    327 => "00111111101000010011110110001100",
    328 => "10111101110011001100110011001101",
    329 => "10111101101111010000001101111011",
    330 => "10111101101111010000001101111011",
    331 => "10111101101111010000001101111011",
    332 => "10111101101111010000001101111011",
    333 => "10111101101111010000001101111011",
    334 => "10111101101111010000001101111011",
    335 => "10111101101111010000001101111011",
    336 => "10111101101111010000001101111011",
    337 => "10111101101111010000001101111011",
    338 => "10111101101111010000001101111011",
    339 => "10111101101111010000001101111011",
    340 => "10111101101111010000001101111011",
    341 => "10111101101111010000001101111011",
    342 => "10111101101111010000001101111011",
    343 => "10111101101111010000001101111011",
    344 => "10111101101111010000001101111011",
    345 => "10111101101111010000001101111011",
    346 => "10111101101111010000001101111011",
    347 => "10111101101111010000001101111011",
    348 => "10111101101111010000001101111011",
    349 => "10111101101111010000001101111011",
    350 => "10111101101111010000001101111011",
    351 => "10111101101111010000001101111011",
    352 => "10111101101111010000001101111011",
    353 => "10111101101111010000001101111011",
    354 => "10111101101111010000001101111011",
    355 => "10111101101111010000001101111011",
    356 => "10111111100000001000110000001100",
    357 => "00111111010010110011100101111001",
    358 => "10111101100101100111100110011111",
    359 => "01000000010001010010001001110110",
    360 => "01000000010001010010001001110110",
    361 => "01000000010001010010001001110110",
    362 => "01000000010001010010001001110110",
    363 => "00111111011001100110011001101000",
    364 => "00111110110101101001101111011100",
    365 => "00111110110101101001101111011100",
    366 => "00111110110101101001101111011100",
    367 => "00111110110101101001101111011100",
    368 => "00111110110101101001101111011100",
    369 => "00111110110101101001101111011100",
    370 => "00111110110101101001101111011100",
    371 => "00111110110101101001101111011100",
    372 => "00111110110101101001101111011100",
    373 => "00111110110101101001101111011100",
    374 => "00111110110101101001101111011100",
    375 => "00111110110101101001101111011100",
    376 => "00111110110101101001101111011100",
    377 => "00111110110101101001101111011100",
    378 => "00111110110101101001101111011100",
    379 => "00111110110101101001101111011100",
    380 => "00111110110101101001101111011100",
    381 => "00111110110101101001101111011100",
    382 => "00111110110101101001101111011100",
    383 => "00111110110101101001101111011100",
    384 => "00111110110101101001101111011100",
    385 => "00111110110101101001101111011100",
    386 => "00111110110101101001101111011100",
    387 => "00111110110101101001101111011100",
    388 => "00111110110101101001101111011100",
    389 => "00111110110101101001101111011100",
    390 => "00111110110101101001101111011100",
    391 => "01000000000111010100000001100100",
    392 => "00111110101001100011100010110001",
    393 => "00111111001110101000011110100001",
    394 => "00111111101000010010011000110100",
    395 => "00111111101000010010011000110100",
    396 => "00111111101000010010011000110100",
    397 => "00111111101000010010011000110100",
    398 => "10111101110011001100110011001101",
    399 => "10111101101111001111001001011001",
    400 => "10111101101111001111001001011001",
    401 => "10111101101111001111001001011001",
    402 => "10111101101111001111001001011001",
    403 => "10111101101111001111001001011001",
    404 => "10111101101111001111001001011001",
    405 => "10111101101111001111001001011001",
    406 => "10111101101111001111001001011001",
    407 => "10111101101111001111001001011001",
    408 => "10111101101111001111001001011001",
    409 => "10111101101111001111001001011001",
    410 => "10111101101111001111001001011001",
    411 => "10111101101111001111001001011001",
    412 => "10111101101111001111001001011001",
    413 => "10111101101111001111001001011001",
    414 => "10111101101111001111001001011001",
    415 => "10111101101111001111001001011001",
    416 => "10111101101111001111001001011001",
    417 => "10111101101111001111001001011001",
    418 => "10111101101111001111001001011001",
    419 => "10111101101111001111001001011001",
    420 => "10111101101111001111001001011001",
    421 => "10111101101111001111001001011001",
    422 => "10111101101111001111001001011001",
    423 => "10111101101111001111001001011001",
    424 => "10111101101111001111001001011001",
    425 => "10111101101111001111001001011001",
    426 => "10111111100000001000101111110100",
    427 => "00111111010010110101011011101100",
    428 => "10111101100101101000000110110101",
    429 => "01000000010001010010000111101010",
    430 => "01000000010001010010000111101010",
    431 => "01000000010001010010000111101010",
    432 => "01000000010001010010000111101010",
    433 => "00111111011001100110011001101000",
    434 => "00111110110101101001110100011000",
    435 => "00111110110101101001110100011000",
    436 => "00111110110101101001110100011000",
    437 => "00111110110101101001110100011000",
    438 => "00111110110101101001110100011000",
    439 => "00111110110101101001110100011000",
    440 => "00111110110101101001110100011000",
    441 => "00111110110101101001110100011000",
    442 => "00111110110101101001110100011000",
    443 => "00111110110101101001110100011000",
    444 => "00111110110101101001110100011000",
    445 => "00111110110101101001110100011000",
    446 => "00111110110101101001110100011000",
    447 => "00111110110101101001110100011000",
    448 => "00111110110101101001110100011000",
    449 => "00111110110101101001110100011000",
    450 => "00111110110101101001110100011000",
    451 => "00111110110101101001110100011000",
    452 => "00111110110101101001110100011000",
    453 => "00111110110101101001110100011000",
    454 => "00111110110101101001110100011000",
    455 => "00111110110101101001110100011000",
    456 => "00111110110101101001110100011000",
    457 => "00111110110101101001110100011000",
    458 => "00111110110101101001110100011000",
    459 => "00111110110101101001110100011000",
    460 => "00111110110101101001110100011000",
    461 => "01000000000111010011111110001010",
    462 => "00111110101001100011100100100110",
    463 => "00111111001110101000011011101101",
    464 => "00111111101000010010011010111000",
    465 => "00111111101000010010011010111000",
    466 => "00111111101000010010011010111000",
    467 => "00111111101000010010011010111000",
    468 => "10111101110011001100110011001101",
    469 => "10111101101111001111001010111011",
    470 => "10111101101111001111001010111011",
    471 => "10111101101111001111001010111011",
    472 => "10111101101111001111001010111011",
    473 => "10111101101111001111001010111011",
    474 => "10111101101111001111001010111011",
    475 => "10111101101111001111001010111011",
    476 => "10111101101111001111001010111011",
    477 => "10111101101111001111001010111011",
    478 => "10111101101111001111001010111011",
    479 => "10111101101111001111001010111011",
    480 => "10111101101111001111001010111011",
    481 => "10111101101111001111001010111011",
    482 => "10111101101111001111001010111011",
    483 => "10111101101111001111001010111011",
    484 => "10111101101111001111001010111011",
    485 => "10111101101111001111001010111011",
    486 => "10111101101111001111001010111011",
    487 => "10111101101111001111001010111011",
    488 => "10111101101111001111001010111011",
    489 => "10111101101111001111001010111011",
    490 => "10111101101111001111001010111011",
    491 => "10111101101111001111001010111011",
    492 => "10111101101111001111001010111011",
    493 => "10111101101111001111001010111011",
    494 => "10111101101111001111001010111011",
    495 => "10111101101111001111001010111011",
    496 => "10111111100000001000101111110100",
    497 => "00111111010010110101011001000110",
    498 => "10111101100101101000000110001000",
    499 => "01000000010001010010000111101110",
    500 => "01000000010001010010000111101110",
    501 => "01000000010001010010000111101110",
    502 => "01000000010001010010000111101110",
    503 => "00111111011001100110011001101000",
    504 => "00111110110101101001110100010100",
    505 => "00111110110101101001110100010100",
    506 => "00111110110101101001110100010100",
    507 => "00111110110101101001110100010100",
    508 => "00111110110101101001110100010100",
    509 => "00111110110101101001110100010100",
    510 => "00111110110101101001110100010100",
    511 => "00111110110101101001110100010100",
    512 => "00111110110101101001110100010100",
    513 => "00111110110101101001110100010100",
    514 => "00111110110101101001110100010100",
    515 => "00111110110101101001110100010100",
    516 => "00111110110101101001110100010100",
    517 => "00111110110101101001110100010100",
    518 => "00111110110101101001110100010100",
    519 => "00111110110101101001110100010100",
    520 => "00111110110101101001110100010100",
    521 => "00111110110101101001110100010100",
    522 => "00111110110101101001110100010100",
    523 => "00111110110101101001110100010100",
    524 => "00111110110101101001110100010100",
    525 => "00111110110101101001110100010100",
    526 => "00111110110101101001110100010100",
    527 => "00111110110101101001110100010100",
    528 => "00111110110101101001110100010100",
    529 => "00111110110101101001110100010100",
    530 => "00111110110101101001110100010100",
    531 => "01000000000111010011111110001100",
    532 => "00111110101001100011100100100011",
    533 => "10111101100101101000000110001000",
    534 => "00111111001110101000011011101101",
    535 => "00111111010011101000101000101010",
    536 => "00111111010011101000101000101010",
    537 => "00000000000000000000000000000000",
    538 => "01000000010010100110001011000100",
    539 => "01000000010010100110001011000100",
    540 => "01000000010010100110001011000100",
    541 => "01000000010010100110001011000100",
    542 => "00111111011001100110011001100110",
    543 => "00111110110010010000111011111000",
    544 => "00111110110010010000111011111000",
    545 => "00111110110010010000111011111000",
    546 => "00111110110010010000111011111000",
    547 => "00111110110010010000111011111000",
    548 => "00111110110010010000111011111000",
    549 => "00111110110010010000111011111000",
    550 => "00111110110010010000111011111000",
    551 => "00111110110010010000111011111000",
    552 => "00111110110010010000111011111000",
    553 => "00111110110010010000111011111000",
    554 => "00111110110010010000111011111000",
    555 => "00111110110010010000111011111000",
    556 => "00111110110010010000111011111000",
    557 => "00111110110010010000111011111000",
    558 => "00111110110010010000111011111000",
    559 => "00111110110010010000111011111000",
    560 => "00111110110010010000111011111000",
    561 => "00111110110010010000111011111000",
    562 => "00111110110010010000111011111000",
    563 => "00111110110010010000111011111000",
    564 => "00111110110010010000111011111000",
    565 => "00111110110010010000111011111000",
    566 => "00111110110010010000111011111000",
    567 => "00111110110010010000111011111000",
    568 => "00111110110010010000111011111000",
    569 => "00111110110010010000111011111000",
    570 => "01000000001001110011111000101010",
    571 => "00111110101000011110100010011011",
    572 => "00111111010000110111000111011101",
    573 => "00111111100110101110010110010110",
    574 => "00111111100110101110010110010110",
    575 => "00111111100110101110010110010110",
    576 => "00111111100110101110010110010110",
    577 => "00111111011001100110011001101000",
    578 => "00111111010000101101111000000011",
    579 => "00111111010000101101111000000011",
    580 => "00111111010000101101111000000011",
    581 => "00111111010000101101111000000011",
    582 => "00111111010000101101111000000011",
    583 => "00111111010000101101111000000011",
    584 => "00111111010000101101111000000011",
    585 => "00111111010000101101111000000011",
    586 => "00111111010000101101111000000011",
    587 => "00111111010000101101111000000011",
    588 => "00111111010000101101111000000011",
    589 => "00111111010000101101111000000011",
    590 => "00111111010000101101111000000011",
    591 => "00111111010000101101111000000011",
    592 => "00111111010000101101111000000011",
    593 => "00111111010000101101111000000011",
    594 => "00111111010000101101111000000011",
    595 => "00111111010000101101111000000011",
    596 => "00111111010000101101111000000011",
    597 => "00111111010000101101111000000011",
    598 => "00111111010000101101111000000011",
    599 => "00111111010000101101111000000011",
    600 => "00111111010000101101111000000011",
    601 => "00111111010000101101111000000011",
    602 => "00111111010000101101111000000011",
    603 => "00111111010000101101111000000011",
    604 => "00111111010000101101111000000011",
    605 => "00111111101110011001000001000110",
    606 => "00111111010100111000110000011011",
    607 => "00111111010111100000101010011001",
    608 => "00111111100010101010011000000110",
    609 => "00111111100010101010011000000110",
    610 => "00111111100010101010011000000110",
    611 => "00111111100010101010011000000110",
    612 => "00111111011001100110011001100110",
    613 => "00111111010000000001110011100001",
    614 => "00111111010000000001110011100001",
    615 => "00111111010000000001110011100001",
    616 => "00111111010000000001110011100001",
    617 => "00111111010000000001110011100001",
    618 => "00111111010000000001110011100001",
    619 => "00111111010000000001110011100001",
    620 => "00111111010000000001110011100001",
    621 => "00111111010000000001110011100001",
    622 => "00111111010000000001110011100001",
    623 => "00111111010000000001110011100001",
    624 => "00111111010000000001110011100001",
    625 => "00111111010000000001110011100001",
    626 => "00111111010000000001110011100001",
    627 => "00111111010000000001110011100001",
    628 => "00111111010000000001110011100001",
    629 => "00111111010000000001110011100001",
    630 => "00111111010000000001110011100001",
    631 => "00111111010000000001110011100001",
    632 => "00111111010000000001110011100001",
    633 => "00111111010000000001110011100001",
    634 => "00111111010000000001110011100001",
    635 => "00111111010000000001110011100001",
    636 => "00111111010000000001110011100001",
    637 => "00111111010000000001110011100001",
    638 => "00111111010000000001110011100001",
    639 => "00111111010000000001110011100001",
    640 => "00111111101011110000001001111000",
    641 => "00111111011011000101011010110101",
    642 => "00111111010111000101110111101110",
    643 => "00111111100010111001001111000010",
    644 => "00111111100010111001001111000010",
    645 => "00111111100010111001001111000010",
    646 => "00111111100010111001001111000010",
    647 => "00111111011001100110011001101000",
    648 => "00111111010000010000011111100000",
    649 => "00111111010000010000011111100000",
    650 => "00111111010000010000011111100000",
    651 => "00111111010000010000011111100000",
    652 => "00111111010000010000011111100000",
    653 => "00111111010000010000011111100000",
    654 => "00111111010000010000011111100000",
    655 => "00111111010000010000011111100000",
    656 => "00111111010000010000011111100000",
    657 => "00111111010000010000011111100000",
    658 => "00111111010000010000011111100000",
    659 => "00111111010000010000011111100000",
    660 => "00111111010000010000011111100000",
    661 => "00111111010000010000011111100000",
    662 => "00111111010000010000011111100000",
    663 => "00111111010000010000011111100000",
    664 => "00111111010000010000011111100000",
    665 => "00111111010000010000011111100000",
    666 => "00111111010000010000011111100000",
    667 => "00111111010000010000011111100000",
    668 => "00111111010000010000011111100000",
    669 => "00111111010000010000011111100000",
    670 => "00111111010000010000011111100000",
    671 => "00111111010000010000011111100000",
    672 => "00111111010000010000011111100000",
    673 => "00111111010000010000011111100000",
    674 => "00111111010000010000011111100000",
    675 => "00111111101011111001100100001100",
    676 => "00111111011010101100010000100110",
    677 => "00111111010111000111101011001000",
    678 => "00111111100010111000001110101100",
    679 => "00111111100010111000001110101100",
    680 => "00111111100010111000001110101100",
    681 => "00111111100010111000001110101100",
    682 => "00111111011001100110011001100110",
    683 => "00111111010000001111100000000101",
    684 => "00111111010000001111100000000101",
    685 => "00111111010000001111100000000101",
    686 => "00111111010000001111100000000101",
    687 => "00111111010000001111100000000101",
    688 => "00111111010000001111100000000101",
    689 => "00111111010000001111100000000101",
    690 => "00111111010000001111100000000101",
    691 => "00111111010000001111100000000101",
    692 => "00111111010000001111100000000101",
    693 => "00111111010000001111100000000101",
    694 => "00111111010000001111100000000101",
    695 => "00111111010000001111100000000101",
    696 => "00111111010000001111100000000101",
    697 => "00111111010000001111100000000101",
    698 => "00111111010000001111100000000101",
    699 => "00111111010000001111100000000101",
    700 => "00111111010000001111100000000101",
    701 => "00111111010000001111100000000101",
    702 => "00111111010000001111100000000101",
    703 => "00111111010000001111100000000101",
    704 => "00111111010000001111100000000101",
    705 => "00111111010000001111100000000101",
    706 => "00111111010000001111100000000101",
    707 => "00111111010000001111100000000101",
    708 => "00111111010000001111100000000101",
    709 => "00111111010000001111100000000101",
    710 => "00111111101011111000111011011010",
    711 => "00111111011010101101111100111100",
    712 => "00111111010111000111100011011111",
    713 => "00111111100010111000010010111100",
    714 => "00111111100010111000010010111100",
    715 => "00111111100010111000010010111100",
    716 => "00111111100010111000010010111100",
    717 => "00111111011001100110011001101000",
    718 => "00111111010000001111100100010011",
    719 => "00111111010000001111100100010011",
    720 => "00111111010000001111100100010011",
    721 => "00111111010000001111100100010011",
    722 => "00111111010000001111100100010011",
    723 => "00111111010000001111100100010011",
    724 => "00111111010000001111100100010011",
    725 => "00111111010000001111100100010011",
    726 => "00111111010000001111100100010011",
    727 => "00111111010000001111100100010011",
    728 => "00111111010000001111100100010011",
    729 => "00111111010000001111100100010011",
    730 => "00111111010000001111100100010011",
    731 => "00111111010000001111100100010011",
    732 => "00111111010000001111100100010011",
    733 => "00111111010000001111100100010011",
    734 => "00111111010000001111100100010011",
    735 => "00111111010000001111100100010011",
    736 => "00111111010000001111100100010011",
    737 => "00111111010000001111100100010011",
    738 => "00111111010000001111100100010011",
    739 => "00111111010000001111100100010011",
    740 => "00111111010000001111100100010011",
    741 => "00111111010000001111100100010011",
    742 => "00111111010000001111100100010011",
    743 => "00111111010000001111100100010011",
    744 => "00111111010000001111100100010011",
    745 => "00111111101011111000111110001000",
    746 => "00111111011010101101110101110001",
    747 => "00111111010111000111100100000001",
    748 => "00111111100010111000010010101010",
    749 => "00111111100010111000010010101010",
    750 => "00111111100010111000010010101010",
    751 => "00111111100010111000010010101010",
    752 => "00111111011001100110011001100110",
    753 => "00111111010000001111100100000000",
    754 => "00111111010000001111100100000000",
    755 => "00111111010000001111100100000000",
    756 => "00111111010000001111100100000000",
    757 => "00111111010000001111100100000000",
    758 => "00111111010000001111100100000000",
    759 => "00111111010000001111100100000000",
    760 => "00111111010000001111100100000000",
    761 => "00111111010000001111100100000000",
    762 => "00111111010000001111100100000000",
    763 => "00111111010000001111100100000000",
    764 => "00111111010000001111100100000000",
    765 => "00111111010000001111100100000000",
    766 => "00111111010000001111100100000000",
    767 => "00111111010000001111100100000000",
    768 => "00111111010000001111100100000000",
    769 => "00111111010000001111100100000000",
    770 => "00111111010000001111100100000000",
    771 => "00111111010000001111100100000000",
    772 => "00111111010000001111100100000000",
    773 => "00111111010000001111100100000000",
    774 => "00111111010000001111100100000000",
    775 => "00111111010000001111100100000000",
    776 => "00111111010000001111100100000000",
    777 => "00111111010000001111100100000000",
    778 => "00111111010000001111100100000000",
    779 => "00111111010000001111100100000000",
    780 => "00111111101011111000111101111100",
    781 => "00111111011010101101110110010000",
    782 => "00111111010111000111100011111110",
    783 => "00111111100010111000010010101100",
    784 => "00111111100010111000010010101100",
    785 => "00111111100010111000010010101100",
    786 => "00111111100010111000010010101100",
    787 => "00111111011001100110011001101000",
    788 => "00111111010000001111100100000011",
    789 => "00111111010000001111100100000011",
    790 => "00111111010000001111100100000011",
    791 => "00111111010000001111100100000011",
    792 => "00111111010000001111100100000011",
    793 => "00111111010000001111100100000011",
    794 => "00111111010000001111100100000011",
    795 => "00111111010000001111100100000011",
    796 => "00111111010000001111100100000011",
    797 => "00111111010000001111100100000011",
    798 => "00111111010000001111100100000011",
    799 => "00111111010000001111100100000011",
    800 => "00111111010000001111100100000011",
    801 => "00111111010000001111100100000011",
    802 => "00111111010000001111100100000011",
    803 => "00111111010000001111100100000011",
    804 => "00111111010000001111100100000011",
    805 => "00111111010000001111100100000011",
    806 => "00111111010000001111100100000011",
    807 => "00111111010000001111100100000011",
    808 => "00111111010000001111100100000011",
    809 => "00111111010000001111100100000011",
    810 => "00111111010000001111100100000011",
    811 => "00111111010000001111100100000011",
    812 => "00111111010000001111100100000011",
    813 => "00111111010000001111100100000011",
    814 => "00111111010000001111100100000011",
    815 => "00111111101011111000111101111110",
    816 => "00111111011010101101110110001101",
    817 => "00111111010111000111100100000001",
    818 => "00111111100010111000010010101010",
    819 => "00111111100010111000010010101010",
    820 => "00111111100010111000010010101010",
    821 => "00111111100010111000010010101010",
    822 => "00111111011001100110011001100110",
    823 => "00111111010000001111100100000000",
    824 => "00111111010000001111100100000000",
    825 => "00111111010000001111100100000000",
    826 => "00111111010000001111100100000000",
    827 => "00111111010000001111100100000000",
    828 => "00111111010000001111100100000000",
    829 => "00111111010000001111100100000000",
    830 => "00111111010000001111100100000000",
    831 => "00111111010000001111100100000000",
    832 => "00111111010000001111100100000000",
    833 => "00111111010000001111100100000000",
    834 => "00111111010000001111100100000000",
    835 => "00111111010000001111100100000000",
    836 => "00111111010000001111100100000000",
    837 => "00111111010000001111100100000000",
    838 => "00111111010000001111100100000000",
    839 => "00111111010000001111100100000000",
    840 => "00111111010000001111100100000000",
    841 => "00111111010000001111100100000000",
    842 => "00111111010000001111100100000000",
    843 => "00111111010000001111100100000000",
    844 => "00111111010000001111100100000000",
    845 => "00111111010000001111100100000000",
    846 => "00111111010000001111100100000000",
    847 => "00111111010000001111100100000000",
    848 => "00111111010000001111100100000000",
    849 => "00111111010000001111100100000000",
    850 => "00111111101011111000111101111100",
    851 => "00111111011010101101110110010000",
    852 => "00111111010111000111100011111110",
    853 => "00111111100010111000010010101100",
    854 => "00111111100010111000010010101100",
    855 => "00111111100010111000010010101100",
    856 => "00111111100010111000010010101100",
    857 => "00111111011001100110011001101000",
    858 => "00111111010000001111100100000011",
    859 => "00111111010000001111100100000011",
    860 => "00111111010000001111100100000011",
    861 => "00111111010000001111100100000011",
    862 => "00111111010000001111100100000011",
    863 => "00111111010000001111100100000011",
    864 => "00111111010000001111100100000011",
    865 => "00111111010000001111100100000011",
    866 => "00111111010000001111100100000011",
    867 => "00111111010000001111100100000011",
    868 => "00111111010000001111100100000011",
    869 => "00111111010000001111100100000011",
    870 => "00111111010000001111100100000011",
    871 => "00111111010000001111100100000011",
    872 => "00111111010000001111100100000011",
    873 => "00111111010000001111100100000011",
    874 => "00111111010000001111100100000011",
    875 => "00111111010000001111100100000011",
    876 => "00111111010000001111100100000011",
    877 => "00111111010000001111100100000011",
    878 => "00111111010000001111100100000011",
    879 => "00111111010000001111100100000011",
    880 => "00111111010000001111100100000011",
    881 => "00111111010000001111100100000011",
    882 => "00111111010000001111100100000011",
    883 => "00111111010000001111100100000011",
    884 => "00111111010000001111100100000011",
    885 => "00111111101011111000111101111110",
    886 => "00111111011010101101110110001101",
    887 => "00111111010111000111100011111110",
    888 => "00111111010111000111100100000001",
    889 => "00111111001000100111001011100000",
    890 => "00111111001000100111001011100000",
    891 => "00111110010011001100110011001101",
    892 => "00000000000000000000000000000000",
    893 => "01000000010010100110001011000100",
    894 => "01000000010010100110001011000100",
    895 => "01000000010010100110001011000100",
    896 => "01000000010010100110001011000100",
    897 => "10111110100110011001100110011000",
    898 => "10111110110010010001000000100010",
    899 => "10111110110010010001000000100010",
    900 => "10111110110010010001000000100010",
    901 => "10111110110010010001000000100010",
    902 => "10111110110010010001000000100010",
    903 => "10111110110010010001000000100010",
    904 => "10111110110010010001000000100010",
    905 => "10111110110010010001000000100010",
    906 => "10111110110010010001000000100010",
    907 => "10111110110010010001000000100010",
    908 => "10111110110010010001000000100010",
    909 => "10111110110010010001000000100010",
    910 => "10111110110010010001000000100010",
    911 => "10111110110010010001000000100010",
    912 => "10111110110010010001000000100010",
    913 => "10111110110010010001000000100010",
    914 => "10111110110010010001000000100010",
    915 => "10111110110010010001000000100010",
    916 => "10111110110010010001000000100010",
    917 => "10111110110010010001000000100010",
    918 => "10111110110010010001000000100010",
    919 => "10111110110010010001000000100010",
    920 => "10111110110010010001000000100010",
    921 => "10111110110010010001000000100010",
    922 => "10111110110010010001000000100010",
    923 => "10111110110010010001000000100010",
    924 => "10111110110010010001000000100010",
    925 => "10111111100010101000101111011100",
    926 => "00111110101000011110100010011011",
    927 => "10111110000001100010000101011011",
    928 => "01000000001110101111101011011110",
    929 => "01000000001110101111101011011110",
    930 => "01000000001110101111101011011110",
    931 => "01000000001110101111101011011110",
    932 => "00111111011001100110011001101000",
    933 => "00111110111010100101011001001100",
    934 => "00111110111010100101011001001100",
    935 => "00111110111010100101011001001100",
    936 => "00111110111010100101011001001100",
    937 => "00111110111010100101011001001100",
    938 => "00111110111010100101011001001100",
    939 => "00111110111010100101011001001100",
    940 => "00111110111010100101011001001100",
    941 => "00111110111010100101011001001100",
    942 => "00111110111010100101011001001100",
    943 => "00111110111010100101011001001100",
    944 => "00111110111010100101011001001100",
    945 => "00111110111010100101011001001100",
    946 => "00111110111010100101011001001100",
    947 => "00111110111010100101011001001100",
    948 => "00111110111010100101011001001100",
    949 => "00111110111010100101011001001100",
    950 => "00111110111010100101011001001100",
    951 => "00111110111010100101011001001100",
    952 => "00111110111010100101011001001100",
    953 => "00111110111010100101011001001100",
    954 => "00111110111010100101011001001100",
    955 => "00111110111010100101011001001100",
    956 => "00111110111010100101011001001100",
    957 => "00111110111010100101011001001100",
    958 => "00111110111010100101011001001100",
    959 => "00111110111010100101011001001100",
    960 => "01000000000100001101011000111100",
    961 => "00111110101011110011111110101111",
    962 => "00111111001100011110010000000101",
    963 => "00111111101001111010100010011000",
    964 => "00111111101001111010100010011000",
    965 => "00111111101001111010100010011000",
    966 => "00111111101001111010100010011000",
    967 => "10111110100110011001100110011000",
    968 => "10111110100100010011000011100110",
    969 => "10111110100100010011000011100110",
    970 => "10111110100100010011000011100110",
    971 => "10111110100100010011000011100110",
    972 => "10111110100100010011000011100110",
    973 => "10111110100100010011000011100110",
    974 => "10111110100100010011000011100110",
    975 => "10111110100100010011000011100110",
    976 => "10111110100100010011000011100110",
    977 => "10111110100100010011000011100110",
    978 => "10111110100100010011000011100110",
    979 => "10111110100100010011000011100110",
    980 => "10111110100100010011000011100110",
    981 => "10111110100100010011000011100110",
    982 => "10111110100100010011000011100110",
    983 => "10111110100100010011000011100110",
    984 => "10111110100100010011000011100110",
    985 => "10111110100100010011000011100110",
    986 => "10111110100100010011000011100110",
    987 => "10111110100100010011000011100110",
    988 => "10111110100100010011000011100110",
    989 => "10111110100100010011000011100110",
    990 => "10111110100100010011000011100110",
    991 => "10111110100100010011000011100110",
    992 => "10111110100100010011000011100110",
    993 => "10111110100100010011000011100110",
    994 => "10111110100100010011000011100110",
    995 => "10111111100001010101001100101100",
    996 => "00111111010000110111000111100100",
    997 => "10111110011000111101010110010001",
    998 => "01000000001001011000010101111000",
    999 => "01000000001001011000010101111000");

  constant ans_lut : lut := (
    0 => "00111111100000000000000000000001",
    1 => "00111110101100101011011111111111",
    2 => "00111110001100101011100000000000",
    3 => "00111101011110011000100011001000",
    4 => "00111100011011100100011011000010",
    5 => "00111011101001100101100001110101",
    6 => "00111010111010000100001000100001",
    7 => "00111010001000100010010011101001",
    8 => "00111001111110101011100010001111",
    9 => "00111001001011110000100010000111",
    10 => "00111000011101000110001101110111",
    11 => "00110111101010101001110011001111",
    12 => "00110110111011100011011101010000",
    13 => "00110110001001100100110110101100",
    14 => "00111101011011100100101011001001",
    15 => "00111100101001100101101101000100",
    16 => "00111011111010000100011000001101",
    17 => "00111011001111101010000000101101",
    18 => "00111010100001010001010001100010",
    19 => "00111001101110011100111110100100",
    20 => "00111001000000011011011111101100",
    21 => "00111000001101010001111000111011",
    22 => "00111000100011110111101001101111",
    23 => "00110111110010000101010010000001",
    24 => "00110111000010111101101010111101",
    25 => "00110110010000110100010100111000",
    26 => "00110101100010000101001001111010",
    27 => "00110100101111100101011010100111",
    28 => "00110100000001001110000100001101",
    29 => "00111111000001100000100111111111",
    30 => "00111110100001100000101000000000",
    31 => "00111110000011000101110011110000",
    32 => "00111100101100101011010100010001",
    33 => "00111100001110110010001110000011",
    34 => "00111011110000111111011111001011",
    35 => "00111011010011010011011010110111",
    36 => "00111010001111000000101001101011",
    37 => "00111001110001001110100110011000",
    38 => "00111001010011100011001111101100",
    39 => "00111000110101111110111001110110",
    40 => "00111000011000100001111010000000",
    41 => "00110111111011001100100110010111",
    42 => "00111101101100101011100000010110",
    43 => "00111101001110110010011010101100",
    44 => "00111100110000111111101100011010",
    45 => "00111011100011101111100000100010",
    46 => "00111011000101011011011011101110",
    47 => "00111010100111001100011100110011",
    48 => "00111010001001000010110011001000",
    49 => "00111001101010111110101110110100",
    50 => "00111000110101110011011110100110",
    51 => "00111000011000010101111100010001",
    52 => "00110111111011000000000100100000",
    53 => "00110111011101110010001110011100",
    54 => "00110111000000010110011001001010",
    55 => "00110110100001111000000100110000",
    56 => "00110110000011011110010111010011",
    57 => "00111110111100001000111011100011",
    58 => "01000010101110111110111110100001",
    59 => "11000010100010001100111001001101",
    60 => "00111111010100000101010101101101",
    61 => "01000011001000101100001010111101",
    62 => "10111110001011110001101111011101",
    63 => "10111110100101111010011011011011",
    64 => "00111111010111110110010111111110",
    65 => "00111110101100101011100110110011",
    66 => "00111110011110011000110110000110",
    67 => "00111100111011100100100100000110",
    68 => "00111100101001100101101110011110",
    69 => "00111100011010000100100011000000",
    70 => "00111100001000100010101100010100",
    71 => "00111010011110101011101011110001",
    72 => "00111010001011110000101111011011",
    73 => "00111001111101000110101001101111",
    74 => "00111001101010101010001101001100",
    75 => "00111001011011100100001010100011",
    76 => "00111001001001100101011100101001",
    77 => "00111111010111110110010111111110",
    78 => "00111101111011100100110100001101",
    79 => "00111101101001100101111001101110",
    80 => "00111101011010000100110010101101",
    81 => "00111011101111101010000111111110",
    82 => "00111011100001010001011011101010",
    83 => "00111011001110011101010011110010",
    84 => "00111011000000011011110011011100",
    85 => "00111010101101010010011011011001",
    86 => "00111001000011110111101111001100",
    87 => "00111000110010000101100001010000",
    88 => "00111000100010111101111010111011",
    89 => "00111000010000110100110010100111",
    90 => "00111000000010000101100011110110",
    91 => "00110111101111100110000110000100",
    92 => "00110111100001001110100111100110",
    93 => "00111110101100101011100110110011",
    94 => "00111110011110011000110110000110",
    95 => "00111100111011100100100100000110",
    96 => "00111100101001100101101110011110",
    97 => "00111100011010000100100011000000",
    98 => "00111100001000100010101100010100",
    99 => "00111010011110101011101011110001",
    100 => "00111010001011110000101111011011",
    101 => "00111001111101000110101001101111",
    102 => "00111001101010101010001101001100",
    103 => "00111001011011100100001010100011",
    104 => "00111001001001100101011100101001",
    105 => "00111110111111000001110010101110",
    106 => "00111101111011100100110100001101",
    107 => "00111101101001100101111001101110",
    108 => "00111101011010000100110010101101",
    109 => "00111011101111101010000111111110",
    110 => "00111011100001010001011011101010",
    111 => "00111011001110011101010011110010",
    112 => "00111011000000011011110011011100",
    113 => "00111010101101010010011011011001",
    114 => "00111001000011110111101111001100",
    115 => "00111000110010000101100001010000",
    116 => "00111000100010111101111010111011",
    117 => "00111000010000110100110010100111",
    118 => "00111000000010000101100011110110",
    119 => "00110111101111100110000110000100",
    120 => "00110111100001001110100111100110",
    121 => "00111110110100111000110110011101",
    122 => "01000100000111000100000000000000",
    123 => "00111010110100011011011100010111",
    124 => "01000100110010000000000000000001",
    125 => "00111010001000111101011100001001",
    126 => "01000101100110010010000000000001",
    127 => "00111001010101011111111011000001",
    128 => "01000100011000010000000000000000",
    129 => "00111010100100011010001010110101",
    130 => "01000100011000010000000000000000",
    131 => "00111010100100011010001010110101",
    132 => "00000000000000000000000000000000",
    133 => "01000000000100000000000000000000",
    134 => "00111111100000000000000000000001",
    135 => "10000000000000000000000000000000",
    136 => "00111111010101010000000101000010",
    137 => "00111111000011100000000011010111",
    138 => "01000100110010000000000000000001",
    139 => "00111010001000111101011100001001",
    140 => "01000100010001000000000000000000",
    141 => "00111010101001110010111100000101",
    142 => "01000100010001000000000000000000",
    143 => "00111010101001110010111100000101",
    144 => "01000011011000010000000000000000",
    145 => "00111011100100011010001010110101",
    146 => "01000011011000010000000000000000",
    147 => "00111011100100011010001010110101",
    148 => "01000011011000010000000000000000",
    149 => "00111011100100011010001010110101",
    150 => "01000100000111000100000000000000",
    151 => "00111010110100011011011100010111",
    152 => "01000100000111000100000000000000",
    153 => "00111010110100011011011100010111",
    154 => "01000100011000010000000000000000",
    155 => "00111010100100011010001010110101",
    156 => "01000100111111010010000000000001",
    157 => "00111010000000010111010000101101",
    158 => "01000101101011111100100000000001",
    159 => "00111001001110100110100111011101",
    160 => "01000100000111000100000000000000",
    161 => "00111010110100011011011100010111",
    162 => "01000010110010000000000000000001",
    163 => "00111100001000111101011100001001",
    164 => "01000010110010000000000000000001",
    165 => "00111100001000111101011100001001",
    166 => "01000100000111000100000000000000",
    167 => "00111010110100011011011100010111",
    168 => "01000011110010000000000000000001",
    169 => "00111011001000111101011100001001",
    170 => "01000011110010000000000000000001",
    171 => "00111011001000111101011100001001",
    172 => "01000011110010000000000000000001",
    173 => "00111011001000111101011100001001",
    174 => "01000011110010000000000000000001",
    175 => "00111011001000111101011100001001",
    176 => "01000011110010000000000000000001",
    177 => "00111011001000111101011100001001",
    178 => "00000000000000000000000000000000",
    179 => "00111111100000000000000000000001",
    180 => "10000000000000000000000000000000",
    181 => "00111111100000000000000000000001",
    182 => "00111111111001100110011001100111",
    183 => "00000000000000000000000000000000",
    184 => "00111101110000000010001000111101",
    185 => "10111110000100110001011000100111",
    186 => "10111111000000100111001000100111",
    187 => "00111111101010010111100010100100",
    188 => "10111110000001100000101011000010",
    189 => "10111100101100101011100100011010",
    190 => "00111011001110110010100011001101",
    191 => "10111001110000111111111001110010",
    192 => "10111010100011101111100011110010",
    193 => "00111001000101011011100010100010",
    194 => "10110111100111001100100111011111",
    195 => "00110110001001000011000010000011",
    196 => "10110100101010111111000010010110",
    197 => "10110111110101110011100011011111",
    198 => "00110110011000010110000110100001",
    199 => "10110100111011000000010100100110",
    200 => "00110011011101110010100100111010",
    201 => "10110010000000010110100111110111",
    202 => "00110000100001111000010111001111",
    203 => "10101111000011011110101101111001",
    204 => "10111101100001100000101011000011",
    205 => "00111100000011000101111010001000",
    206 => "10111011101100101011011000010101",
    207 => "00111010001110110010010110100011",
    208 => "10111000110000111111101100100001",
    209 => "00110111010011010011101101011111",
    210 => "10111001001111000000101101111100",
    211 => "00110111110001001110101111010100",
    212 => "10110110010011100011011101101111",
    213 => "00110100110101111111001101011101",
    214 => "10110011011000100010010011101100",
    215 => "00110001111011001101000110101001",
    216 => "10111110000001101101000000011011",
    217 => "10111101001010101000011010111111",
    218 => "00111010111000110010111001111001",
    219 => "00111101101111100111110101101111",
    220 => "10111110000101000110011110101011",
    221 => "10111111000000100101110100000000",
    222 => "00111111101010000010011010100001",
    223 => "00111111100101011001101111100110",
    224 => "00111110010011011100111111001001",
    225 => "00111101101001010111011001101111",
    226 => "00111100100010010011001011110000",
    227 => "00111011110111001001101001001011",
    228 => "00111011001100010101101010011011",
    229 => "00111010100011101001010110000001",
    230 => "00111010000100000101110101010001",
    231 => "00111001011010000001111111001100",
    232 => "00111000101110101001110111011101",
    233 => "00111000000101100000011111100001",
    234 => "00110111011100010011110000101001",
    235 => "00110110110000011111000011111001",
    236 => "00111101100010010011010101000010",
    237 => "00111100110111001001111000000110",
    238 => "00111100001100010101110110011011",
    239 => "00111011010110111000011000001110",
    240 => "00111010101100000111110010000110",
    241 => "00111010000011011110001011110110",
    242 => "00111001011001000010001111010001",
    243 => "00111000101101110110100111011001",
    244 => "00111000101001010011101010010111",
    245 => "00111000000001001101011000000110",
    246 => "00110111010101011001011001100111",
    247 => "00110110101010111011011011001100",
    248 => "00110110000010100000110011000000",
    249 => "00110101010111011111100010000100",
    250 => "00110100101100100111010000101011",
    251 => "01000000000101101000101101010010",
    252 => "00111111010000000001000101110111",
    253 => "00111111000100000001101000110100",
    254 => "00111101000101010011111110011000",
    255 => "10111110000000010100101010110010",
    256 => "10111110001101001100110110101100",
    257 => "00111111011011000101100000010001",
    258 => "10111101101110100000000101011000",
    259 => "10111100011110000000000111101011",
    260 => "00111010101101000011001010110010",
    261 => "10111001000000101110110111000111",
    262 => "10111010010001100110010111001110",
    263 => "00111000100100000010011100000010",
    264 => "10110110110100010111101000110010",
    265 => "00110101000110000011001111100010",
    266 => "10110011010111010010110011111110",
    267 => "10110111100101010101001111110111",
    268 => "00110101110110001111111110010100",
    269 => "10110100000111011010101011010101",
    270 => "00110010011001010001110111100110",
    271 => "10110000101001100111100011101101",
    272 => "00101110111100011110100101111000",
    273 => "10101101001011111100010011100110",
    274 => "10111101001110100000000101011001",
    275 => "00111011100001110010010111110100",
    276 => "10111011011101111111110110111011",
    277 => "00111001101101000010111110100111",
    278 => "10111000000000101110101110010001",
    279 => "00110110001111100011111110101111",
    280 => "10111001000000100111100010110101",
    281 => "00110111001111011001100011000110",
    282 => "10110101100010011100000111111111",
    283 => "00110011110010000010111101011001",
    284 => "10110010000100010111001101110011",
    285 => "00110000010100110101110101001010",
    286 => "10111101101110101000010010110101",
    287 => "10111101100101111101110001011011",
    288 => "00111011101101000010101101100010",
    289 => "00111101101110110000111101011000",
    290 => "10111110000101110000001101001011",
    291 => "10111111000000100000010111110000",
    292 => "00111111101001011010010110001001",
    293 => "00111111100100110101101011101010",
    294 => "00111110010101101101001110111001",
    295 => "00111101101101000100011010100111",
    296 => "00111100100011110011010101110111",
    297 => "00111011111100000101101001000011",
    298 => "00111011010010011011001000111011",
    299 => "00111010101010010100000111001100",
    300 => "00111010000101101011000000110010",
    301 => "00111001011111001110011111010011",
    302 => "00111000110101000011101011110011",
    303 => "00111000001100100001100011001100",
    304 => "00110111100101010111010000000101",
    305 => "00110110111110101101010100101100",
    306 => "00111101100011110011011111100011",
    307 => "00111100111100000101111001010011",
    308 => "00111100010010011011010110100100",
    309 => "00111011011001010010001111000010",
    310 => "00111010110000000100100101100101",
    311 => "00111010001000010101110001100001",
    312 => "00111001100001110110100010101100",
    313 => "00111000111000110100001011111001",
    314 => "00111000101011000111011101110001",
    315 => "00111000000100001011101001111011",
    316 => "00110111011100101110011100101001",
    317 => "00110110110010111101011000011111",
    318 => "00110110001010110000110110010010",
    319 => "00110101100011111000101011001111",
    320 => "00110100111100001110100110000000",
    321 => "01000000000011110111100101011101",
    322 => "00111111001110100110011110001000",
    323 => "00111111000001111011101010011011",
    324 => "00111101000110010001001010010111",
    325 => "10111110000000110110011001111010",
    326 => "10111110001111000001011110011100",
    327 => "00111111011100000001101010111101",
    328 => "10111101101111010000001101111011",
    329 => "10111100011111000000010011000101",
    330 => "00111010101110100001001011110010",
    331 => "10111001000010010110001010000100",
    332 => "10111010010010011001101101000000",
    333 => "00111000100101001101101001011100",
    334 => "10110110110110111100111001111000",
    335 => "00110101001000100100101001101011",
    336 => "10110011011011111010011001001100",
    337 => "10110111100101111011111000111110",
    338 => "00110101111000000001001100001000",
    339 => "10110100001001010111000100011001",
    340 => "00110010011101000100110101111111",
    341 => "10110000101101000110000010001001",
    342 => "00101111000001010010110110111001",
    343 => "10101101010001001010100100100010",
    344 => "10111101001111010000001101111100",
    345 => "00111011100010111000111000100100",
    346 => "10111011011111000000000010000011",
    347 => "00111001101110100000111111001110",
    348 => "10111000000010010110000000110010",
    349 => "00110110010010101101101111000110",
    350 => "10111001000001001001010011101010",
    351 => "00110111010000111100011101111101",
    352 => "10110101100100001000110011110001",
    353 => "00110011110101010111010000001010",
    354 => "10110010000111011001100110010010",
    355 => "00110000011010001011100100001011",
    356 => "10111101101111011000110101010011",
    357 => "10111101100101100111100110011111",
    358 => "00111011101100001110010110000000",
    359 => "00111101101110110010011000001000",
    360 => "10111110000101101111001010101011",
    361 => "10111111000000100000100011101000",
    362 => "00111111101001011011010100001110",
    363 => "00111111100100110110100011100001",
    364 => "00111110010101101001101111011101",
    365 => "00111101101100111110100011110011",
    366 => "00111100100011110001000000111011",
    367 => "00111011111011111101110101010110",
    368 => "00111011010010010001010100001111",
    369 => "00111010101010001001001000000111",
    370 => "00111010000101101000100100000011",
    371 => "00111001011111000110010001011110",
    372 => "00111000110100111001010110010000",
    373 => "00111000001100010101111111010111",
    374 => "00110111100101001011001000011011",
    375 => "00110110111110010100111011010101",
    376 => "00111101100011110001001010100101",
    377 => "00111100111011111110000101100010",
    378 => "00111100010010010001100001110011",
    379 => "00111011011001001110100000101101",
    380 => "00111010101111111110010101110011",
    381 => "00111010001000001101111010100011",
    382 => "00111001100001101101110000001101",
    383 => "00111000111000100001110000011100",
    384 => "00111000101011000100101010011001",
    385 => "00111000000100000110111101000001",
    386 => "00110111011100100010100111100000",
    387 => "00110110110010110000001001110001",
    388 => "00110110001010100010111110100011",
    389 => "00110101100011101010101101101111",
    390 => "00110100111011110011010001010111",
    391 => "01000000000011111010001101111010",
    392 => "00111111001110101000011110100001",
    393 => "00111111000001111110100101011110",
    394 => "00111101000110001111110001101110",
    395 => "10111110000000110101101001101110",
    396 => "10111110001110111110110100110111",
    397 => "00111111011100000000010101010010",
    398 => "10111101101111001111001001011001",
    399 => "10111100011110111110110111101101",
    400 => "00111010101110011111000100111000",
    401 => "10111001000010010011110100101100",
    402 => "10111010010010011000100011111010",
    403 => "00111000100101001011111101100001",
    404 => "10110110110110111001001010111000",
    405 => "00110101001000100000111110011100",
    406 => "10110011011011110011100111000011",
    407 => "10110111100101111011000001111101",
    408 => "00110101110111111110101001101011",
    409 => "10110100001001010100010000100000",
    410 => "00110010011100111111010011110111",
    411 => "10110000101101000000111011011000",
    412 => "00101111000001001110010101011011",
    413 => "10101101010001000010110001111100",
    414 => "10111101001111001111001001011010",
    415 => "00111011100010110111010011011001",
    416 => "10111011011110111110100110101100",
    417 => "00111001101110011110111000010101",
    418 => "10111000000010010011101011011011",
    419 => "00110110010010101001001001000101",
    420 => "10111001000001001000100011100101",
    421 => "00110111010000111010010000000000",
    422 => "10110101100100000110010110100101",
    423 => "00110011110101010010011010101111",
    424 => "10110010000111010101001000110001",
    425 => "00110000011010000011101010010101",
    426 => "10111101101111010111110000001110",
    427 => "10111101100101101000000110110101",
    428 => "00111011101100001111100010000100",
    429 => "00111101101110110010010110000011",
    430 => "10111110000101101111001100001100",
    431 => "10111111000000100000100011010101",
    432 => "00111111101001011011010010110110",
    433 => "00111111100100110110100010010010",
    434 => "00111110010101101001110100011001",
    435 => "00111101101100111110101100000101",
    436 => "00111100100011110001000100001101",
    437 => "00111011111011111110000000010111",
    438 => "00111011010010010001100010000110",
    439 => "00111010101010001001010111100111",
    440 => "00111010000101101000100111100001",
    441 => "00111001011111000110011101000110",
    442 => "00111000110100111001100100110111",
    443 => "00111000001100010110001111101101",
    444 => "00110111100101001011011001100011",
    445 => "00110110111110010101011101110001",
    446 => "00111101100011110001001101111000",
    447 => "00111100111011111110010000100101",
    448 => "00111100010010010001101111101100",
    449 => "00111011011001001110100101111110",
    450 => "00111010101111111110011110101000",
    451 => "00111010001000001110000101101001",
    452 => "00111001100001101101111100100111",
    453 => "00111000111000100010001010011100",
    454 => "00111000101011000100101110010110",
    455 => "00111000000100000111000011101010",
    456 => "00110111011100100010111000001101",
    457 => "00110110110010110000011100011011",
    458 => "00110110001010100011010010000111",
    459 => "00110101100011101011000001011011",
    460 => "00110100111011110011110111111000",
    461 => "01000000000011111010001010001011",
    462 => "00111111001110101000011011101101",
    463 => "00111111000001111110100001010111",
    464 => "00111101000110001111110011101011",
    465 => "10111110000000110101101010110010",
    466 => "10111110001110111110111000100110",
    467 => "00111111011100000000010111001100",
    468 => "10111101101111001111001010111011",
    469 => "10111100011110111110111001110000",
    470 => "00111010101110011111000111111010",
    471 => "10111001000010010011111000000010",
    472 => "10111010010010011000100101100010",
    473 => "00111000100101001011111111111011",
    474 => "10110110110110111001010000001101",
    475 => "00110101001000100001000011101100",
    476 => "10110011011011110011110000110000",
    477 => "10110111100101111011000011001011",
    478 => "00110101110111111110101101010010",
    479 => "10110100001001010100010100100000",
    480 => "00110010011100111111011011101111",
    481 => "10110000101101000001000010101001",
    482 => "00101111000001001110011011110111",
    483 => "10101101010001000010111101000010",
    484 => "10111101001111001111001010111100",
    485 => "00111011100010110111010101101001",
    486 => "10111011011110111110101000101110",
    487 => "00111001101110011110111011010101",
    488 => "10111000000010010011101110110000",
    489 => "00110110010010101001001111101000",
    490 => "10111001000001001000100100101010",
    491 => "00110111010000111010010011001011",
    492 => "10110101100100000110011010000110",
    493 => "00110011110101010010100001101010",
    494 => "10110010000111010101001111001010",
    495 => "00110000011010000011110101101001",
    496 => "10111101101111010111110001110000",
    497 => "10111101100101101000000110001000",
    498 => "00111011101100001111100000011010",
    499 => "00111101101110110010010110000111",
    500 => "10111110000101101111001100001001",
    501 => "10111111000000100000100011010110",
    502 => "00111111101001011011010010110111",
    503 => "00111111100100110110100010010011",
    504 => "00111110010101101001110100010101",
    505 => "00111101101100111110101011111110",
    506 => "00111100100011110001000100001010",
    507 => "00111011111011111110000000001110",
    508 => "00111011010010010001100001111011",
    509 => "00111010101010001001010111011010",
    510 => "00111010000101101000100111011110",
    511 => "00111001011111000110011100111100",
    512 => "00111000110100111001100100101011",
    513 => "00111000001100010110001111011111",
    514 => "00110111100101001011011001010100",
    515 => "00110110111110010101011101010011",
    516 => "00111101100011110001001101110101",
    517 => "00111100111011111110010000011100",
    518 => "00111100010010010001101111100001",
    519 => "00111011011001001110100101111001",
    520 => "00111010101111111110011110100000",
    521 => "00111010001000001110000101100000",
    522 => "00111001100001101101111100011101",
    523 => "00111000111000100010001010000111",
    524 => "00111000101011000100101110010011",
    525 => "00111000000100000111000011100101",
    526 => "00110111011100100010111000000000",
    527 => "00110110110010110000011100001101",
    528 => "00110110001010100011010001111000",
    529 => "00110101100011101011000001001011",
    530 => "00110100111011110011110111011000",
    531 => "01000000000011111010001010001101",
    532 => "00111111001110101000011011101101",
    533 => "00111011101100001111100000011010",
    534 => "00111111000001111110100001010111",
    535 => "10111101011100101101101011101100",
    536 => "00111111000101100111110100111110",
    537 => "00000000000000000000000000000000",
    538 => "00111101110000000010001000111101",
    539 => "10111110000100110001011000100111",
    540 => "10111111000000100111001000100111",
    541 => "00111111101010010111100010100100",
    542 => "00111111100101101100110000011010",
    543 => "00111110010010010000111011111001",
    544 => "00111101100111011110100010000011",
    545 => "00111100100001100000011111001000",
    546 => "00111011110100101000011111100101",
    547 => "00111011001001010101100100000010",
    548 => "00111010100000011101110010001101",
    549 => "00111010000011010000011111001011",
    550 => "00111001010111011000011010111011",
    551 => "00111000101011011111101110111101",
    552 => "00111000000010001010010011010100",
    553 => "00110111010101101010001011010000",
    554 => "00110110101010001001001001100010",
    555 => "00111101100001100000101000001100",
    556 => "00111100110100101000101101110100",
    557 => "00111100001001010101101111001101",
    558 => "00111011010101100111010000101100",
    559 => "00111010101010000110110111000000",
    560 => "00111010000001000100100000000101",
    561 => "00111001010011111100100010010000",
    562 => "00111000101000110011000010011111",
    563 => "00111000101000010110100110110111",
    564 => "00110111111111011000101011100010",
    565 => "00110111010001110010000011011111",
    566 => "00110110100111000110010001110100",
    567 => "00110101111101011010100000001000",
    568 => "00110101010000001110111101001011",
    569 => "00110100100101111000011100101010",
    570 => "01000000000110101000001100111110",
    571 => "00111111010000110111000111011101",
    572 => "00111111000101010011011010101001",
    573 => "00111101000100110000110011100101",
    574 => "10111110000000000000110101111001",
    575 => "10111110001100001010010000100000",
    576 => "00111111011010100001111101011011",
    577 => "00111111010011110100000110101101",
    578 => "00111110110000101101111000000100",
    579 => "00111110100101000101010100111110",
    580 => "00111101000000011110011100110110",
    581 => "00111100110001011100001110111110",
    582 => "00111100100101101000100111011000",
    583 => "00111100011001010010111000000110",
    584 => "00111010100010001011000000001011",
    585 => "00111010010100000001011111100101",
    586 => "00111010000111100110011010010010",
    587 => "00111001111100010010011000110011",
    588 => "00111001101101111001000000010100",
    589 => "00111001100010111011101001100000",
    590 => "00111110000000011110100101101000",
    591 => "00111101110001011100011100010101",
    592 => "00111101100101101000110001100011",
    593 => "00111011110011111101100110011111",
    594 => "00111011100111100011011100101011",
    595 => "00111011011100001101111000001000",
    596 => "00111011001101110101100100100101",
    597 => "00111011000010111001000010001111",
    598 => "00111001000111000111000101001001",
    599 => "00111000111011100010101100001011",
    600 => "00111000101101010100101100101010",
    601 => "00111000100010100000000000101111",
    602 => "00111000010100100001011110100011",
    603 => "00111000000111111110110000011100",
    604 => "00110111111100110111011100111100",
    605 => "00111111100001100101100110000001",
    606 => "00111111010111100000101010011001",
    607 => "00111111010000001001011001100010",
    608 => "00111101000000111010000000001001",
    609 => "10111101111011011001100000111101",
    610 => "10111110000101000001011000101110",
    611 => "00111111010110010100101111001111",
    612 => "00111111010000000001110011100001",
    613 => "00111110000000000001001101010001",
    614 => "00111101110000000011100111011111",
    615 => "00111101100100000100000100010110",
    616 => "00111011110011001110100110000010",
    617 => "00111011100110011100011000111111",
    618 => "00111011011001101100110000010000",
    619 => "00111011001011010011001100010101",
    620 => "00111011000000011111100111011001",
    621 => "00111001000110100011101100110010",
    622 => "00111000111001110111101110010111",
    623 => "00111000101011011011011011001110",
    624 => "00111000100000100101110010110011",
    625 => "00111000010000111010100001110110",
    626 => "00111000000100101101010001101011",
    627 => "00110111110111000101111111000001",
    628 => "00111110110000000001110011100010",
    629 => "00111110100100000010101101010101",
    630 => "00111101000000000001000100100111",
    631 => "00111100110000000011011010100000",
    632 => "00111100100100000011111010100111",
    633 => "00111100010110000111111010000110",
    634 => "00111010100001101100000101101111",
    635 => "00111010010010100100000010001110",
    636 => "00111010000101111100011100111011",
    637 => "00111001111000111100110100010111",
    638 => "00111001101010101111001110000100",
    639 => "00111001100000000100100111101100",
    640 => "00111111011011101011001100010011",
    641 => "00111111010111000101110111101110",
    642 => "00111111001111011011000110010011",
    643 => "00111101000001001000000110111011",
    644 => "10111101111011101011010010010011",
    645 => "10111110000101011010111100100000",
    646 => "00111111010110100101000011101001",
    647 => "00111111010000010000011111100000",
    648 => "00111110000000001010111111111011",
    649 => "00111101110000100001000101000011",
    650 => "00111101100100100101010011111100",
    651 => "00111011110011011110010000101001",
    652 => "00111011100110110011111101011000",
    653 => "00111011011010100001111100010000",
    654 => "00111011001100001000100010011110",
    655 => "00111011000001010001110001101101",
    656 => "00111001000110101111011111011010",
    657 => "00111000111010011011001100111111",
    658 => "00111000101100000011011101010011",
    659 => "00111000100001001101111100100001",
    660 => "00111000010010000110000010011100",
    661 => "00111000000101110001011011111111",
    662 => "00110111111000111101100111111000",
    663 => "00111110110000010000011111100001",
    664 => "00111110100100011000110011100000",
    665 => "00111101000000001010110111001111",
    666 => "00111100110000100000110111111101",
    667 => "00111100100100100101001010000011",
    668 => "00111100010111001010100101101010",
    669 => "00111010100001110110011001000101",
    670 => "00111010010011000011000010001001",
    671 => "00111010000110011111011011011111",
    672 => "00111001111010000010111110110101",
    673 => "00111001101011110001001100011011",
    674 => "00111001100001000000001011001010",
    675 => "00111111011100000110101111010110",
    676 => "00111111010111000111101011001000",
    677 => "00111111001111011110001101000010",
    678 => "00111101000001000111001001110101",
    679 => "10111101111011101010000101100100",
    680 => "10111110000101011001001101101011",
    681 => "00111111010110100011111101001100",
    682 => "00111111010000001111100000000101",
    683 => "00111110000000001010010101101001",
    684 => "00111101110000011111000101100011",
    685 => "00111101100100100011000011110000",
    686 => "00111011110011011101001101000000",
    687 => "00111011100110110010010111011001",
    688 => "00111011011010011110010101100101",
    689 => "00111011001100000100111010100110",
    690 => "00111011000001001110010111001100",
    691 => "00111001000110101110101100100000",
    692 => "00111000111010011000110011011110",
    693 => "00111000101100000000101111101011",
    694 => "00111000100001001011001101111111",
    695 => "00111000010010000000111001100000",
    696 => "00111000000101101100110010011010",
    697 => "00110111111000110101011100011001",
    698 => "00111110110000001111100000000110",
    699 => "00111110100100010111010011111001",
    700 => "00111101000000001010001100111101",
    701 => "00111100110000011110111000011101",
    702 => "00111100100100100010111001111000",
    703 => "00111100010111000110000011110100",
    704 => "00111010100001110101101100100110",
    705 => "00111010010011000000111011111111",
    706 => "00111010000110011101000011110010",
    707 => "00111001111001111110001101110110",
    708 => "00111001101011101100101101000001",
    709 => "00111001100000111100000111001001",
    710 => "00111111011100000100111000001000",
    711 => "00111111010111000111100011011111",
    712 => "00111111001111011101111111111000",
    713 => "00111101000001000111001101110111",
    714 => "10111101111011101010001010101000",
    715 => "10111110000101011001010100111111",
    716 => "00111111010110100100000001110110",
    717 => "00111111010000001111100100010011",
    718 => "00111110000000001010011000011101",
    719 => "00111101110000011111001110000010",
    720 => "00111101100100100011001101010110",
    721 => "00111011110011011101010001100000",
    722 => "00111011100110110010011110001011",
    723 => "00111011011010011110100100111011",
    724 => "00111011001100000101001010000001",
    725 => "00111011000001001110100101101110",
    726 => "00111001000110101110101111111001",
    727 => "00111000111010011000111101101100",
    728 => "00111000101100000000111011001111",
    729 => "00111000100001001011011001100111",
    730 => "00111000010010000001001111011001",
    731 => "00111000000101101101000110001101",
    732 => "00110111111000110101111111001110",
    733 => "00111110110000001111100100010100",
    734 => "00111110100100010111011010010000",
    735 => "00111101000000001010001111110001",
    736 => "00111100110000011111000000111100",
    737 => "00111100100100100011000011011110",
    738 => "00111100010111000110010111000110",
    739 => "00111010100001110101101111100011",
    740 => "00111010010011000001000100111010",
    741 => "00111010000110011101001101110111",
    742 => "00111001111001111110100010000111",
    743 => "00111001101011101101000000001000",
    744 => "00111001100000111100011000011011",
    745 => "00111111011100000101000000000010",
    746 => "00111111010111000111100100000001",
    747 => "00111111001111011110000000110011",
    748 => "00111101000001000111001101100110",
    749 => "10111101111011101010001010010011",
    750 => "10111110000101011001010100100000",
    751 => "00111111010110100100000001100011",
    752 => "00111111010000001111100100000000",
    753 => "00111110000000001010011000010001",
    754 => "00111101110000011111001101011101",
    755 => "00111101100100100011001100101011",
    756 => "00111011110011011101010001001100",
    757 => "00111011100110110010011101101100",
    758 => "00111011011010011110100011110101",
    759 => "00111011001100000101001000111011",
    760 => "00111011000001001110100100101100",
    761 => "00111001000110101110101111101001",
    762 => "00111000111010011000111100111101",
    763 => "00111000101100000000111010011010",
    764 => "00111000100001001011011000110010",
    765 => "00111000010010000001001101110110",
    766 => "00111000000101101101000100110011",
    767 => "00110111111000110101111100110000",
    768 => "00111110110000001111100100000001",
    769 => "00111110100100010111011001110011",
    770 => "00111101000000001010001111100100",
    771 => "00111100110000011111000000010101",
    772 => "00111100100100100011000010110010",
    773 => "00111100010111000110010101101110",
    774 => "00111010100001110101101111010110",
    775 => "00111010010011000001000100010010",
    776 => "00111010000110011101001101001010",
    777 => "00111001111001111110100000101100",
    778 => "00111001101011101100111110110010",
    779 => "00111001100000111100010111001101",
    780 => "00111111011100000100111111011111",
    781 => "00111111010111000111100011111110",
    782 => "00111111001111011110000000101101",
    783 => "00111101000001000111001101101000",
    784 => "10111101111011101010001010010101",
    785 => "10111110000101011001010100100100",
    786 => "00111111010110100100000001100101",
    787 => "00111111010000001111100100000011",
    788 => "00111110000000001010011000010011",
    789 => "00111101110000011111001101100011",
    790 => "00111101100100100011001100110010",
    791 => "00111011110011011101010001001111",
    792 => "00111011100110110010011101110001",
    793 => "00111011011010011110100100000000",
    794 => "00111011001100000101001001000110",
    795 => "00111011000001001110100100110110",
    796 => "00111001000110101110101111101100",
    797 => "00111000111010011000111101000101",
    798 => "00111000101100000000111010100011",
    799 => "00111000100001001011011000111010",
    800 => "00111000010010000001001110000101",
    801 => "00111000000101101101000101000001",
    802 => "00110111111000110101111101001000",
    803 => "00111110110000001111100100000100",
    804 => "00111110100100010111011001110111",
    805 => "00111101000000001010001111100110",
    806 => "00111100110000011111000000011011",
    807 => "00111100100100100011000010111001",
    808 => "00111100010111000110010101111100",
    809 => "00111010100001110101101111011000",
    810 => "00111010010011000001000100011000",
    811 => "00111010000110011101001101010001",
    812 => "00111001111001111110100000111010",
    813 => "00111001101011101100111110111111",
    814 => "00111001100000111100010111011001",
    815 => "00111111011100000100111111100110",
    816 => "00111111010111000111100100000001",
    817 => "00111111001111011110000000110011",
    818 => "00111101000001000111001101100110",
    819 => "10111101111011101010001010010011",
    820 => "10111110000101011001010100100000",
    821 => "00111111010110100100000001100011",
    822 => "00111111010000001111100100000000",
    823 => "00111110000000001010011000010001",
    824 => "00111101110000011111001101011101",
    825 => "00111101100100100011001100101011",
    826 => "00111011110011011101010001001100",
    827 => "00111011100110110010011101101100",
    828 => "00111011011010011110100011110101",
    829 => "00111011001100000101001000111011",
    830 => "00111011000001001110100100101100",
    831 => "00111001000110101110101111101001",
    832 => "00111000111010011000111100111101",
    833 => "00111000101100000000111010011010",
    834 => "00111000100001001011011000110010",
    835 => "00111000010010000001001101110110",
    836 => "00111000000101101101000100110011",
    837 => "00110111111000110101111100110000",
    838 => "00111110110000001111100100000001",
    839 => "00111110100100010111011001110011",
    840 => "00111101000000001010001111100100",
    841 => "00111100110000011111000000010101",
    842 => "00111100100100100011000010110010",
    843 => "00111100010111000110010101101110",
    844 => "00111010100001110101101111010110",
    845 => "00111010010011000001000100010010",
    846 => "00111010000110011101001101001010",
    847 => "00111001111001111110100000101100",
    848 => "00111001101011101100111110110010",
    849 => "00111001100000111100010111001101",
    850 => "00111111011100000100111111011111",
    851 => "00111111010111000111100011111110",
    852 => "00111111001111011110000000101101",
    853 => "00111101000001000111001101101000",
    854 => "10111101111011101010001010010101",
    855 => "10111110000101011001010100100100",
    856 => "00111111010110100100000001100101",
    857 => "00111111010000001111100100000011",
    858 => "00111110000000001010011000010011",
    859 => "00111101110000011111001101100011",
    860 => "00111101100100100011001100110010",
    861 => "00111011110011011101010001001111",
    862 => "00111011100110110010011101110001",
    863 => "00111011011010011110100100000000",
    864 => "00111011001100000101001001000110",
    865 => "00111011000001001110100100110110",
    866 => "00111001000110101110101111101100",
    867 => "00111000111010011000111101000101",
    868 => "00111000101100000000111010100011",
    869 => "00111000100001001011011000111010",
    870 => "00111000010010000001001110000101",
    871 => "00111000000101101101000101000001",
    872 => "00110111111000110101111101001000",
    873 => "00111110110000001111100100000100",
    874 => "00111110100100010111011001110111",
    875 => "00111101000000001010001111100110",
    876 => "00111100110000011111000000011011",
    877 => "00111100100100100011000010111001",
    878 => "00111100010111000110010101111100",
    879 => "00111010100001110101101111011000",
    880 => "00111010010011000001000100011000",
    881 => "00111010000110011101001101010001",
    882 => "00111001111001111110100000111010",
    883 => "00111001101011101100111110111111",
    884 => "00111001100000111100010111011001",
    885 => "00111111011100000100111111100110",
    886 => "00111111010111000111100100000001",
    887 => "00111111001111011110000000101101",
    888 => "00111111001111011110000000110011",
    889 => "00111111000010111110011101111111",
    890 => "00111111000010111110011110000001",
    891 => "00111111000110011001100110011010",
    892 => "00000000000000000000000000000000",
    893 => "00111101110000000010001000111101",
    894 => "10111110000100110001011000100111",
    895 => "10111111000000100111001000100111",
    896 => "00111111101010010111100010100100",
    897 => "10111110110010010001000000100010",
    898 => "10111101100001100000101011010011",
    899 => "00111100110100101000110111100101",
    900 => "10111100001001010101111010101101",
    901 => "10111011010101100111010101101010",
    902 => "00111010101010000110111110110100",
    903 => "10111010000001000100101001010010",
    904 => "00111001010011111100110101100010",
    905 => "10111000101000110011010101011010",
    906 => "10111000101000010110101010100110",
    907 => "00110111111111011000110111010001",
    908 => "10110111010001110010010001010011",
    909 => "00110110100111000110100000010010",
    910 => "10110101111101011010111100100011",
    911 => "00110101010000001111010111111110",
    912 => "10110100100101111000110101001101",
    913 => "10111110010010010001000000100011",
    914 => "00111101100111011110101001010111",
    915 => "10111100100001100000100010001111",
    916 => "00111011110100101000101001010110",
    917 => "10111011001001010101101111100010",
    918 => "00111010100000011101111110010000",
    919 => "10111010000011010000100010011100",
    920 => "00111001010111011000100101001100",
    921 => "10111000101011011111111011000011",
    922 => "00111000000010001010011111111110",
    923 => "10110111010101101010100100000110",
    924 => "00110110101010001001100000111101",
    925 => "10111110110101000001010000100000",
    926 => "10111110000001100010000101011011",
    927 => "00111100100011001000110111100000",
    928 => "00111101101100011000001000011111",
    929 => "10111110000111010100000100110101",
    930 => "10111110111111111110001011001010",
    931 => "00111111101000000011101000101000",
    932 => "00111111100011100111101001000101",
    933 => "00111110011010100101011001001101",
    934 => "00111101110101101000000111100001",
    935 => "00111100100111000011011011111001",
    936 => "00111100000011101111111011101000",
    937 => "00111011100000101110010100110100",
    938 => "00111010111011111010001101000011",
    939 => "00111010001001000101111110010111",
    940 => "00111001100101100111011011001001",
    941 => "00111001000010011011101101001100",
    942 => "00111000011111000010011101000010",
    943 => "00110111111001101101000011100010",
    944 => "00110111010100110100100010111101",
    945 => "00111101100111000011100110011100",
    946 => "00111101000011110000000101010010",
    947 => "00111100100000101110011101101010",
    948 => "00111011011110011111001100011000",
    949 => "00111010111001001100110001110110",
    950 => "00111010010100010111000000000100",
    951 => "00111001101111111011011011111101",
    952 => "00111001001011110111110111100011",
    953 => "00111000101111000010000100101011",
    954 => "00111000001011000011010110111100",
    955 => "00110111100111011010001100101011",
    956 => "00110111000100000100110001001001",
    957 => "00110110100001000001011001011111",
    958 => "00110101111100011101000111110011",
    959 => "00110101010111010101101101101100",
    960 => "01000000000000011110110111111101",
    961 => "00111111001100011110010000000101",
    962 => "00111110111101110011101000110100",
    963 => "00111101000111110010101001101000",
    964 => "10111110000001101010001010101110",
    965 => "10111110010001111101000100010110",
    966 => "00111111011101011101001010001111",
    967 => "10111110100100010011000011100110",
    968 => "10111101010000011001011010100010",
    969 => "00111100010110111001011010011000",
    970 => "10111011011110010001010001111100",
    971 => "10111011000110101101110100111110",
    972 => "00111010001011111010100111001010",
    973 => "10111001010001110100000101110010",
    974 => "00111000011000100000010001000010",
    975 => "10110111100000000010111110010101",
    976 => "10111000011010010001111110010010",
    977 => "00110111100001000011011101101001",
    978 => "10110110100101011111100101001000",
    979 => "00110101101010100001110110101111",
    980 => "10110100110000001111011010011101",
    981 => "00110011110110101110000100010101",
    982 => "10110010111110000100011010011000",
    983 => "10111110000100010011000011100111",
    984 => "00111101001001001011000011011101",
    985 => "10111100010000011001001101011101",
    986 => "00111011010110111001001011100011",
    987 => "10111010011110010001000001000111",
    988 => "00111001100011010100000111001011",
    989 => "10111001110010111010111110000001",
    990 => "00111000111001110000101010100000",
    991 => "10111000000000110000100100100110",
    992 => "00110111000101001010001001101100",
    993 => "10110110001010001001100011000111",
    994 => "00110101001111110011110101111010",
    995 => "10111110100101010011011001011010",
    996 => "10111110011000111101010110010001",
    997 => "00111101010010101100010001110001",
    998 => "00111101100111010010001011111111",
    999 => "10111110001001011000110011111110");

  component fmul is
    port (A : in std_logic_vector (31 downto 0);
          B : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          C : out std_logic_vector (31 downto 0));
  end component fmul;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal s_b : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (4 downto 0) of std_logic_vector (31 downto 0);
  signal cc : buff := (others => (others => '0'));
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
  signal i_isRunning : std_logic := '0';
  signal i_result : std_logic := '1';
begin  -- architecture fmul_tb

  i_fmul : fmul port map (s_a,s_b,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk) is
    variable ss : character;
    variable count : integer := 4;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      case state is
        when "00" =>
          state <= "01";
        when "01" =>
          state <= "11";
        when "11" =>
          state <= "10";
        when others =>
          state <= "00";
      end case;
      s_a <= a_lut (addr);
      s_b <= b_lut (addr);
      cc(conv_integer(state)) <= ans_lut (addr);      
      if i_isRunning = '1' then  -- rising clock edge
        ccc <= cc (conv_integer (state));
        if (ccc = c or state /= "00") and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 5 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;
  end process ram_loop;

end architecture;
