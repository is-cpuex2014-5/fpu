library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity fsqrt_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity fsqrt_tb;

architecture testbench of fsqrt_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "00110001011110111010101111011000",
    1 => "01101010110111011000001000001011",
    2 => "01101001111111110111001100100000",
    3 => "00011111111101000000110111100001",
    4 => "00011111100110110001111110100101",
    5 => "00101111111111011100000011111100",
    6 => "01110100111111100101100101010100",
    7 => "01101111101111111110010001000101",
    8 => "00110101111110111010110100101100",
    9 => "01100111111111110101010110111101",
    10 => "01110101101111100101100011011011",
    11 => "00011011110111111110111010101011",
    12 => "01001111111111111000010001001000",
    13 => "01111110110111110010011111011111",
    14 => "01101100110101101010100100101001",
    15 => "01110010111011111111110000101010",
    16 => "00110011111111111011010011111000",
    17 => "01110100110011110010000011010111",
    18 => "01101000100001110000110110101100",
    19 => "00111101100111101001001100011111",
    20 => "00111100110111010111110101011111",
    21 => "01111101101110011001101001100010",
    22 => "01010011110101110010001011011111",
    23 => "01101101101110110011111011100011",
    24 => "00001101101111010010111101101100",
    25 => "01101111011111011011000001001011",
    26 => "01110110110001110100000110010011",
    27 => "00100100011010111000110011111000",
    28 => "01111101101011010100100110100011",
    29 => "00010111111111111010011100010010",
    30 => "01110111010111110110010000000100",
    31 => "01011111101111010100111101110011",
    32 => "01011111011101101010110000001001",
    33 => "00001011111111100010111101101111",
    34 => "01011010011011111110001000010100",
    35 => "01011111101011110100111011011010",
    36 => "00100011111111110011000001001000",
    37 => "01000111111110111000011001101001",
    38 => "00110100110110110100001101001000",
    39 => "00111001011111111100001000101111",
    40 => "00110001111100100100001001000100",
    41 => "00111101011101110110101100101001",
    42 => "01110110010111001000101100011101",
    43 => "00011111100111111101110101110111",
    44 => "00111000101001110100111100010000",
    45 => "01101111111010110100101011010100",
    46 => "01100110011111110100000100101100",
    47 => "01101101111111110001101000001000",
    48 => "00111111010111101111101010101110",
    49 => "01101100010111110101010110110101",
    50 => "01011100011110110001010011101101",
    51 => "01111100111110110000001000101100",
    52 => "01011001011111000100011110110100",
    53 => "00110011111111111110001110010100",
    54 => "00101110111111001010100010101010",
    55 => "00001111011101110100000000010001",
    56 => "00111011111111111010010001110010",
    57 => "00011101111110110110011011010110",
    58 => "00110101111011000000110001111001",
    59 => "00111011111101111011110100000101",
    60 => "01011111000111110001000001101110",
    61 => "00001111101111111101010110010110",
    62 => "01111101011011001011001101101110",
    63 => "01101111011101110010100100000101",
    64 => "00111111111111110000100011001100",
    65 => "00111010101111110101011011100110",
    66 => "01110110111111111000010100110101",
    67 => "01110111001111110111101011010010",
    68 => "01111001011010010101011111100111",
    69 => "01011111111010101000110011010101",
    70 => "01111110001110011000010011001001",
    71 => "01011001010111101101000010010111",
    72 => "01011100110111100111010111101000",
    73 => "01011011011110011010101100111101",
    74 => "00111101111010101001101111010101",
    75 => "00111011111100111101010001000000",
    76 => "01011111111001011010101001001001",
    77 => "01101001111111111101101001001011",
    78 => "00000111110110011011101010010011",
    79 => "01111011111111011010000101101111",
    80 => "01111101111011110100011001000000",
    81 => "01101011101111111000111111110000",
    82 => "00111100111101110110101101101010",
    83 => "01011001000110010101000111110000",
    84 => "00111011011010111010001011000100",
    85 => "01110011110101101000100111010000",
    86 => "01111101111111101010001110010000",
    87 => "00110011101101101100000010011010",
    88 => "01101110001101101101000000111101",
    89 => "01001111111111110011110001110010",
    90 => "00011111111111001001100101001000",
    91 => "01111101110111111101010100001111",
    92 => "01111001110101011000111111000100",
    93 => "00111011100111010110101110010101",
    94 => "00110100111110011110100110100110",
    95 => "01010111111110110100001111011000",
    96 => "01000101001111100010010100011010",
    97 => "01101100111001110110011010100010",
    98 => "01010111101101110001001100101000",
    99 => "01110111111101111110010101000001",
    100 => "00011011101001010011100100000111",
    101 => "00011101110111111001011101011011",
    102 => "00111111101110100011010000010100",
    103 => "01011001101111100101101101111110",
    104 => "01100001111110001110101110110000",
    105 => "00100100111101110010001011100110",
    106 => "00011111100011110101110010111001",
    107 => "00011111101111111010101011110101",
    108 => "01010011111100111110110111110110",
    109 => "00111111011001011101111110011000",
    110 => "01011101111111111110001110101100",
    111 => "01110111110010010001100100111000",
    112 => "01111101111101110010100010100111",
    113 => "01111011101110110111000011101111",
    114 => "01110111110001110011011011011000",
    115 => "01111101111111011110000010100111",
    116 => "01110110111000000000010110111100",
    117 => "00111011011111111110101001101011",
    118 => "01101011111011011101000000111111",
    119 => "01111111010111101010010100100110",
    120 => "00111111011111111110110001111000",
    121 => "00111001111111110010110001000010",
    122 => "00001111111011011111110010101011",
    123 => "01011111111101111010010100100001",
    124 => "01110111011100111001001100110001",
    125 => "01111011100011111011100000110100",
    126 => "01111110101111110100101000010001",
    127 => "00111101010100000111010011110011",
    128 => "01101010101100110110101001111001",
    129 => "01110111011111111101011110010110",
    130 => "01011010010000100111100010101100",
    131 => "01111100111010111100011010111010",
    132 => "01110100110110110101111100111011",
    133 => "00101000111011110100110111011011",
    134 => "01111101111111110000101100111010",
    135 => "01110111100111101001001111100011",
    136 => "01111110111111110110011000101101",
    137 => "00111011101101111000110111001101",
    138 => "01110110110001100010110101000010",
    139 => "01011111110111110000010101100000",
    140 => "01110111111111011000110001101010",
    141 => "01101111111110111010110000010101",
    142 => "00010111010110111100101100101101",
    143 => "01101101111100011001100011011010",
    144 => "00100101111101001011101000101111",
    145 => "01000111101111110000011101011101",
    146 => "00111000111000010101110101111111",
    147 => "00001011110111100010100111110000",
    148 => "01111011111000010001101111010110",
    149 => "01111110111011110000001111010111",
    150 => "00010111111111110010110100001011",
    151 => "00101101011111111111001001000100",
    152 => "01101111110110100101101010000000",
    153 => "01111111011111011111001101100010",
    154 => "01011101100111111011100010111010",
    155 => "00111111111111111011010010010010",
    156 => "01011111101111010110000111011100",
    157 => "01101111111101111100001101000010",
    158 => "00011010111011001000011010101011",
    159 => "01010101110111010010101111101001",
    160 => "01111011111111111011010011110101",
    161 => "01101110110110110000000100111000",
    162 => "01111111011111111010011011001100",
    163 => "01011111101101111010011101011010",
    164 => "01111110111101110011010010111001",
    165 => "01110111100111110110111000011000",
    166 => "01101111010101000011011100110010",
    167 => "01101110011010110111110100110010",
    168 => "00111111111111110110001111101011",
    169 => "01110111111111100010010110001100",
    170 => "01101110111110100110000110111010",
    171 => "01111111001111110010100100111101",
    172 => "01101101010111010101001001101111",
    173 => "01010101100111010000100011000011",
    174 => "01110110110111111110110001000110",
    175 => "00100011111110100101100000100101",
    176 => "01111110101111110110101110000011",
    177 => "00111011111111111111100101010101",
    178 => "00101111001111110010101000010101",
    179 => "01111101011101010010101100101111",
    180 => "00101101111110110011001010111011",
    181 => "01011011101111010001100001111111",
    182 => "00101101111101111000101010110000",
    183 => "01101110101111101010010110100110",
    184 => "01100111011111111010100000111100",
    185 => "01101110110111111001011010000000",
    186 => "01101101001000011101011001110010",
    187 => "01111100101111111010101001010100",
    188 => "01111101111111000111001011001000",
    189 => "00111110111111001100011110011001",
    190 => "00011111111111101110101111000101",
    191 => "00101111111111111100100110000000",
    192 => "01111011111111100001000110010100",
    193 => "00111011001101111111101000101000",
    194 => "00011110111010011001000000111000",
    195 => "01110111110111111100101100111100",
    196 => "01011111011100111001111111001111",
    197 => "01110110110101010111011101010001",
    198 => "01000110111101110111000100000110",
    199 => "00111110111110001110011100000111",
    200 => "00111010111111011111001011010001",
    201 => "00111111101011110000010110001110",
    202 => "01010101000011110001000101000000",
    203 => "01101100101111010110010001100010",
    204 => "01011001110111010001110010000101",
    205 => "01101001111111110001100111010011",
    206 => "00101010110111111100010110101111",
    207 => "01101010011011101101000010010100",
    208 => "01101001111101110111110100101001",
    209 => "01111011111111000000111001010101",
    210 => "00011111110101111100111011110000",
    211 => "01110111010111110101000100001011",
    212 => "01011101011010111001010001001011",
    213 => "01111010101111110111110010111001",
    214 => "01010110111010110011001111010010",
    215 => "00101111111011001111101000011111",
    216 => "01111110110110111100011100001001",
    217 => "00001111111111111111111010111001",
    218 => "01001111001111100001100100111001",
    219 => "00111011011011111011000010111110",
    220 => "01011111111101010111110111100101",
    221 => "01111011110111110000000111000010",
    222 => "00101111011001101011001110110010",
    223 => "00111100101111110000010100010001",
    224 => "01101111111111100010101110101111",
    225 => "00110110111100111111100011100000",
    226 => "01111101111111110001000000101101",
    227 => "01111111001001101001000100010110",
    228 => "00101110111111111000011011001000",
    229 => "00011111110101111010011100001100",
    230 => "01100111111011101110000011001110",
    231 => "01001111011111111010011000110001",
    232 => "00111110100001100100001101000010",
    233 => "01111110111010110000100011110111",
    234 => "01101010111101100000111001110010",
    235 => "00111101010010111001110011100111",
    236 => "01001101111100110000100000001001",
    237 => "01101011111010001101010000011100",
    238 => "00010111110111111100110010001100",
    239 => "01110110011110111100001010000111",
    240 => "01111011101110010101101100111101",
    241 => "00110101011011110110111100111001",
    242 => "01111101101011111000100010010101",
    243 => "01011110111100111001110101111101",
    244 => "00011101111110111011000000001010",
    245 => "01011100111101111011001111000110",
    246 => "00001111011110110101011010100101",
    247 => "01101111111101110000011010010111",
    248 => "01011011110111000111010011111011",
    249 => "00111110000101110010011110011001",
    250 => "01111001000111011101000100000100",
    251 => "00011111111101110100101000000010",
    252 => "00111011111110111100001111011000",
    253 => "01101111001100101000001101100100",
    254 => "01111101101111011100010111100001",
    255 => "01101111111111101111100100101010",
    256 => "01010110111100110110000011111010",
    257 => "01111101111101111101000110010001",
    258 => "00111111010101110001001001110000",
    259 => "01110011111011110100110001101000",
    260 => "01111010011101011011010101111000",
    261 => "00111111010111110110111010001001",
    262 => "01000111111111110010110010111000",
    263 => "00011001101100111000100011111101",
    264 => "00111110101110011011011101100000",
    265 => "01100101011111100011101010110110",
    266 => "01111111011110101010010001010010",
    267 => "01011101111110110010101101110111",
    268 => "01111010010110001000100101000000",
    269 => "01011001010110100010101100101111",
    270 => "00000111010110110010101100001101",
    271 => "01101111111110110100000001101101",
    272 => "00111111111111111001001111001001",
    273 => "00101111111011100011011111101100",
    274 => "00111011111111111111111001110111",
    275 => "01111110110010011011101011011011",
    276 => "01101101110110111111110010010100",
    277 => "00101111111110111100010100001010",
    278 => "01110101111110110010001101101101",
    279 => "01111110010101101100101111100001",
    280 => "01111011111111110000010110101110",
    281 => "01010011010111111011110100000111",
    282 => "01111101110100101011010111111101",
    283 => "00111111001001110111101100011100",
    284 => "00110111011111110110000111010000",
    285 => "01110101111111111111100000100001",
    286 => "00101111111111101110010111000110",
    287 => "00111101001000010000110100100010",
    288 => "01111011111111111100010010010101",
    289 => "01101101111110011001100100100101",
    290 => "01110110011111110100011111100000",
    291 => "01011111101011010111100110110000",
    292 => "00111111111111110000100010111110",
    293 => "01011011101111111101100100111001",
    294 => "01011111011101111111100101010011",
    295 => "01011011001011001000010011000011",
    296 => "01111011111100011001000100011001",
    297 => "01000111111010011010100001110001",
    298 => "01111101011111111011000100001100",
    299 => "01001111101011011111111000010001",
    300 => "00111110110011111001101011111000",
    301 => "00101111110101010111110001011011",
    302 => "01110110101111111111100000011001",
    303 => "01010111111101010010010110101001",
    304 => "01111110111110111001001000110100",
    305 => "01111011101110010100100011011001",
    306 => "01011111111011100010110101111011",
    307 => "01111100101110100100110110111001",
    308 => "01010101110111111111100000000011",
    309 => "01111011101100010001011100100110",
    310 => "00111100111011111110010000001001",
    311 => "01110111110111111101000010110101",
    312 => "01111110101111110010010110100011",
    313 => "01101110011111111010010100000001",
    314 => "01111010011111101011010101100110",
    315 => "01111011011111111001101011110000",
    316 => "01011011011001110100100011110010",
    317 => "01110011110110111000010001010000",
    318 => "01101011111110111101010000000111",
    319 => "00111001111101111000001101110100",
    320 => "01100000111111010011100011011101",
    321 => "00001101111000110101001010110100",
    322 => "00111000010110110110111001101011",
    323 => "00001011110110111000001001100001",
    324 => "00111111111111110000101100111010",
    325 => "01110111001111111001110001001110",
    326 => "01100011100111111000011111011111",
    327 => "01111011111111101011010001000101",
    328 => "01110011001011111000100011110111",
    329 => "00110011111011110000000010100011",
    330 => "01101101100011111101011000010111",
    331 => "01111001101111001100111000011111",
    332 => "01101101111011101001101010000001",
    333 => "01101111100111110010010011000011",
    334 => "01111111011111110010110101011101",
    335 => "01101111111101100000000101010100",
    336 => "01110111101111110011111111111110",
    337 => "01101111010111110010010011011001",
    338 => "01110111110111011000110010000110",
    339 => "00011101110110010000100100100100",
    340 => "01011111100101111001011011100100",
    341 => "01111101110111111110111110111001",
    342 => "01011001111010101101000010111000",
    343 => "01101111011001011001101110010000",
    344 => "00001011101001100111100100011101",
    345 => "01101101111110100110101010100010",
    346 => "00111111101111110111111001110111",
    347 => "01111011111111110001011111111011",
    348 => "01111001000111111000001100010011",
    349 => "01111100111111110001000011101010",
    350 => "01111101111111011001011101010001",
    351 => "00111011111010010001101001110011",
    352 => "01110101011110110111111010001100",
    353 => "01011101111110111001001111001110",
    354 => "01110110011110110110100000110111",
    355 => "01111111011111001100110011101001",
    356 => "01111110111111110010110101000101",
    357 => "01011001110110100101101101110000",
    358 => "01101100011111110000000111111100",
    359 => "01011010110110011100110000101111",
    360 => "01111101100111111100001010110000",
    361 => "01010110111111111001001001001000",
    362 => "01010111101011110111100111000100",
    363 => "01111101111110100011001101001100",
    364 => "01110111110101101111011000101110",
    365 => "01011001111101000100000000111100",
    366 => "01011111001011101111110000110010",
    367 => "01111011111110110010101010100111",
    368 => "01011111111111110001100011000001",
    369 => "01101101111110111010001000010101",
    370 => "01111011010011101111101101000011",
    371 => "01100010111111111101111101101100",
    372 => "01110111111111101111101111011000",
    373 => "00101100111110111100110011001100",
    374 => "00111011111101100011111010111101",
    375 => "00001001111101011111001110010111",
    376 => "00011111011111101011100101100011",
    377 => "01011011111110110101111011010000",
    378 => "01001101000111110101101101000010",
    379 => "01011011001011101100001010110110",
    380 => "00111111111111010101110000100111",
    381 => "00110111111110110111001001100100",
    382 => "01101111011110110111011111000110",
    383 => "01101111111101100000101011011010",
    384 => "01110010111111111000010011010000",
    385 => "01111101110100110010101100011000",
    386 => "01111110111011101001010000111110",
    387 => "01111100000110111000111110010001",
    388 => "01110110111101100100110100111111",
    389 => "00001011101011010110110100011110",
    390 => "01111101111011011000011101100001",
    391 => "01111110101110001000000010001100",
    392 => "00011110110011100100001001110110",
    393 => "01101101101111111110011010111100",
    394 => "01110111011111110000010100110000",
    395 => "00001111111011111100100000100111",
    396 => "01010111011101110011010011011001",
    397 => "01101111111110011000001000010101",
    398 => "01100111111001101101101001101100",
    399 => "01111001110110110110011001000110",
    400 => "01111011110101110100011110011001",
    401 => "01111111001110111110111111000111",
    402 => "00101111110011111111111000100010",
    403 => "00100110110010111010001111001010",
    404 => "00101111111111111010010010010000",
    405 => "01111110111101011100001100001001",
    406 => "01010100111011110000010101101010",
    407 => "00010111111011100110111011111110",
    408 => "00110110111111111001101110101001",
    409 => "00111111111100111100010100101010",
    410 => "01101111111111110100101100100000",
    411 => "01011000111111110011001111110101",
    412 => "00101110101010101011000000100011",
    413 => "01111011110011100000110110111001",
    414 => "01101111101111010001011110000010",
    415 => "01111000111111111000101000001000",
    416 => "00100101111110100000010011100011",
    417 => "01011100110011010110011111000111",
    418 => "01111001100001111001110011101100",
    419 => "01110111010001110101001110000001",
    420 => "01101011111101101110100010110001",
    421 => "01010011111111110110111101110000",
    422 => "00101111111111011101011101110110",
    423 => "01100101111111111001111000111000",
    424 => "01100010111111111000011100110001",
    425 => "01010111110110101011011011001110",
    426 => "01011111101110101011110101110011",
    427 => "01111011110111101001010011000101",
    428 => "01111111000110110100011110000110",
    429 => "01110011110111111000010101010011",
    430 => "01101110001111110010100111000100",
    431 => "01111011101110100101110010000101",
    432 => "01111011111111100010110011100011",
    433 => "01001101101111110110010011010110",
    434 => "01110111111011001110001011011010",
    435 => "00111110111111110110111101000111",
    436 => "00110111111111100101110001111111",
    437 => "00110111111110110111101010001110",
    438 => "01110101101110100101100011011010",
    439 => "01111101111111011010011110110000",
    440 => "01101101111101110111000000010011",
    441 => "00110111111111111000010001101010",
    442 => "01100111111101001010101000101111",
    443 => "01111101111101100110100111001010",
    444 => "01100011110010110110110001011011",
    445 => "01110111010111111011000100110101",
    446 => "01111111011101110000101000010010",
    447 => "01110111110111010111101110011110",
    448 => "00101100011101110011001010110000",
    449 => "01111011011110110000011111001001",
    450 => "00111111111011010000110111011100",
    451 => "00101110010111011111010011111110",
    452 => "00111111111101011100100010010000",
    453 => "01011100011110110111101101010101",
    454 => "00011110110111000111011111010111",
    455 => "00111111111111010000101001011110",
    456 => "01011110111011010100111111110010",
    457 => "01111011111001110001001110001100",
    458 => "01110011011111111010111111000111",
    459 => "01111010011001110001010000101000",
    460 => "01111111010011011000111111100110",
    461 => "01110111001101101000101010010001",
    462 => "01111101110111111110110111100011",
    463 => "01110001110011111100000110100010",
    464 => "01111111011101110110100100110011",
    465 => "01000111111010110001111110100000",
    466 => "01111010011010010011110110001011",
    467 => "01011111111101010110010000101000",
    468 => "01101001101111110010100000011011",
    469 => "01101111111111111000110100101111",
    470 => "01111011100110111001011011010100",
    471 => "01111010011111110111000100111000",
    472 => "00010111011110011010110000011110",
    473 => "00111101110101010010111001000000",
    474 => "01111110111111110010001100101010",
    475 => "01100101101111010000101001110010",
    476 => "01100111111111010011010000110110",
    477 => "01111011100111010001110001101010",
    478 => "00001011111011111101110010010100",
    479 => "01111011101011110100100000001101",
    480 => "01111100111101010110011100101000",
    481 => "01110011011111101010001101000000",
    482 => "01101111011100010101011000110100",
    483 => "01011110111111111101110100010011",
    484 => "00011101101111100001000100011000",
    485 => "00100110111111110101101001100001",
    486 => "01110011010110001011110000001110",
    487 => "01001111111111110011111000010101",
    488 => "00111110011111110110001101101101",
    489 => "01111011110110101000100111101011",
    490 => "01111110111111110010101011111001",
    491 => "01110111100100111000100101001100",
    492 => "01110111111111110111100011000010",
    493 => "01111111001101100011111010001100",
    494 => "01111110101111110110011110011111",
    495 => "00101001111110110000101000111101",
    496 => "01011000111111100001100110111101",
    497 => "00111011110101110011001101100011",
    498 => "00111100011111110101101000100101",
    499 => "00011011101111011101010001100110",
    500 => "01011101111110110010000001101000",
    501 => "01001111110111110111110010101100",
    502 => "01111110101111111000000010000111",
    503 => "00010111101101110101011010001110",
    504 => "00111011010110110010001000100010",
    505 => "00011111101101111010011101111011",
    506 => "01111011101011111101010010011011",
    507 => "00101111111100010000010010110100",
    508 => "00111101011101111010110100001100",
    509 => "01111111010001111011010001000101",
    510 => "01110110111100010000101011000000",
    511 => "01000010110110110001011110010001",
    512 => "01111110111011100011100101111100",
    513 => "00011111001111101010111101001111",
    514 => "00011011010011010011101100011100",
    515 => "00111111110101111110001011011110",
    516 => "01101111101011111001110011111001",
    517 => "01110100111111000011110111010000",
    518 => "01011011011011110001010010110001",
    519 => "01011111111011111011110100000001",
    520 => "01111110100011110100000100101100",
    521 => "00111011110101110100110110011000",
    522 => "00111011011101110000010100111001",
    523 => "01111110110011111110101001101111",
    524 => "00110101111011111101010001110111",
    525 => "01101111111111101111100011011111",
    526 => "01111110111111011110101110011111",
    527 => "00101111011111011111111011100000",
    528 => "00010011110101111010001011100001",
    529 => "01111101110101110010110011111000",
    530 => "01111101101110111011010111000011",
    531 => "01111011111111010010111101011001",
    532 => "01100011111100010101111111000000",
    533 => "01111001110111111000001111100101",
    534 => "00111111111101110000000011001101",
    535 => "01110011110010110010000010101110",
    536 => "01101011011010110011010100011010",
    537 => "01100010110100100010001101110001",
    538 => "00111111011010101101110010100010",
    539 => "01100101111111111001110100000011",
    540 => "00111110001111011101000000101101",
    541 => "01001110111010110100110111001100",
    542 => "01111101010010010000101010111000",
    543 => "01111101011000010000110011001100",
    544 => "01111111011111101110111001100110",
    545 => "00011111111111110000100101011100",
    546 => "01101111111010111101011110010111",
    547 => "01100001010101001111100000000000",
    548 => "01011101111111010000110010010100",
    549 => "00110111011111110110101111011110",
    550 => "01111011111111110110111000010101",
    551 => "01111100011111000100010010101101",
    552 => "01011011110011110001011110010111",
    553 => "01010101111111000110101111101011",
    554 => "00110111010101011111100111100000",
    555 => "00110111011111111111010011100000",
    556 => "01100011111111110110100100100001",
    557 => "01111110111011111101100101101001",
    558 => "01101110001111111111011000000011",
    559 => "00001111101110100001011010111101",
    560 => "01101011111110111110000100100010",
    561 => "01110111101111111101001000110110",
    562 => "00101011101110101101001010001011",
    563 => "00111111100110110101001010111011",
    564 => "01101111111111100101111100111001",
    565 => "01111101111101110111110000101101",
    566 => "00111111100111110101011001011001",
    567 => "01100011111111100011100001011101",
    568 => "01110111111110100010110101000101",
    569 => "01111110111101111000010000100100",
    570 => "01111001110101101110101101111111",
    571 => "00011010101010110010011110010011",
    572 => "01100111110111110110001101101001",
    573 => "01111101000111110111010111110101",
    574 => "01001111100101010001101101100001",
    575 => "01011101101001101101110101101011",
    576 => "01101011100111111010111101100111",
    577 => "00011111111110110101011100001101",
    578 => "01100110101011000011000100001011",
    579 => "01110111111111100100111100110100",
    580 => "01010100110011011101111010101111",
    581 => "00110011010111010101011101011011",
    582 => "01111011111101010001011010011100",
    583 => "00010111010111110000101111010001",
    584 => "01011111010110100100100001111101",
    585 => "00100111111011001100110101011100",
    586 => "01111110111010111000111110111110",
    587 => "00101100011011110010111110110101",
    588 => "01101110111001110010100001011100",
    589 => "01100111111110110010000001101001",
    590 => "01110111100111110111110111110101",
    591 => "00011111100100000100101001100011",
    592 => "01011101010011010101010110101100",
    593 => "01101110111110101100101011001100",
    594 => "00011101011101111111000110000011",
    595 => "00011011110111111010111110001010",
    596 => "01111001111011000110001110101010",
    597 => "01111110110010110011001011111010",
    598 => "01111110110011001111100000001110",
    599 => "01100101111011111101111100101100",
    600 => "01111101011111100001101011111110",
    601 => "01100101101111111100010010011100",
    602 => "01111011011111010001101001000001",
    603 => "01101101100001100011111101101100",
    604 => "01011111011111100100010101011010",
    605 => "01100111110011101110111010110100",
    606 => "00111101111011110101001111000000",
    607 => "01111110101110110110000000110110",
    608 => "01110111101010001000110101110110",
    609 => "00111011101111101000001110010101",
    610 => "01101011011101011011001111100100",
    611 => "01110111111111110000001001011010",
    612 => "01010111110111110100100011001000",
    613 => "01101100111101111100011001111110",
    614 => "00100110101111100011111110001000",
    615 => "01111101111011111011110110101000",
    616 => "00011010111110100100000100111000",
    617 => "01011111101100011111000101111010",
    618 => "01111101101101011110010011000100",
    619 => "01110010111001110110110101101110",
    620 => "00011010111111111110100001101101",
    621 => "00101011111111110010101110010111",
    622 => "01011111111110110011000101111001",
    623 => "01110111100011011101011011111010",
    624 => "00111010111011111100110110101010",
    625 => "01011111111011110110110010010111",
    626 => "00001001111011111100110011100000",
    627 => "01110110110111111000111001111100",
    628 => "01110011101101001110000011011101",
    629 => "00111111111110110011011000111010",
    630 => "01111110101111100100110101000001",
    631 => "00111101011110110110111110101010",
    632 => "01111110111111001011011101111010",
    633 => "00111011111010110100011111100101",
    634 => "01111110110100101100101100101111",
    635 => "01001101111011111010011100000111",
    636 => "01101010010111110001011011000001",
    637 => "01000010111111110011010101000100",
    638 => "01111010111111110011100100100001",
    639 => "00011110011101100011100010001101",
    640 => "01111111001111111111011001011101",
    641 => "01110010111111101111000110011010",
    642 => "01110111111011110100101100000000",
    643 => "01110101111010010110100100011110",
    644 => "01111011011111110001000000001110",
    645 => "01111101010100100011010110000111",
    646 => "01010010101110111011110010010100",
    647 => "00011111110111011000000101110010",
    648 => "00011101111111111001001010001011",
    649 => "01100111110111110010011011011001",
    650 => "00110111111101111000110111111000",
    651 => "01100100101111110111110000111010",
    652 => "00111111001000110011001000100111",
    653 => "01100110111110110000100111010101",
    654 => "00111011111101100000100001011001",
    655 => "01111010110101011111000001101101",
    656 => "01011110111111110111001010011001",
    657 => "01110110000000011010110010101110",
    658 => "01110101110101111100111100000000",
    659 => "01111100111111111011000011110000",
    660 => "01001011111110111111011000001101",
    661 => "01011101111111111100011011110000",
    662 => "00101110011110110011010010100001",
    663 => "00111110111011111111110110100101",
    664 => "01000111010010110010100101001111",
    665 => "00011111011110111101010110101011",
    666 => "00111110101010010000010101000100",
    667 => "01011111011001110011110010110011",
    668 => "00110011101000111101111101110111",
    669 => "01100011110111011100101101011111",
    670 => "00101001100010101000011100010001",
    671 => "01111101111000110010111000100110",
    672 => "00000011101111111001101001010000",
    673 => "01111101101111001110111000110111",
    674 => "01110101101101101011100110111010",
    675 => "00111111010001011000010100011010",
    676 => "01111110101110110110010110110110",
    677 => "00110100000111110001101000000101",
    678 => "01101111101011111000101001111110",
    679 => "00101111111111110100101100100010",
    680 => "00111011110111010111101111111101",
    681 => "00111111101111111010100000010011",
    682 => "01111111011110111011101011010010",
    683 => "01111111010011111000111110111101",
    684 => "01111110111011101000011011110101",
    685 => "01111111011101010110011011110011",
    686 => "00111101111000110101010011111110",
    687 => "01010111111111111110010000100010",
    688 => "01011111111111110001000010000010",
    689 => "01001111100111010100110001000100",
    690 => "01111111001101111011011111011100",
    691 => "01101111101111101110111010110010",
    692 => "01111001111110110111100001110011",
    693 => "00111011000110000000110001100000",
    694 => "01011111100111110101000010101100",
    695 => "01110111011110001001001111010000",
    696 => "01110101011110110010000101100100",
    697 => "01001101101111110110111101000011",
    698 => "01011101110110111000011011111000",
    699 => "00111111101010110001101011000101",
    700 => "01001111111010110111001010111011",
    701 => "00011011100011111100001111100001",
    702 => "01001010111110111001100110100101",
    703 => "00101111010111101110001001010100",
    704 => "01111011111111111011000101101110",
    705 => "00111101011011110110011000010111",
    706 => "01111011111101010110101101000100",
    707 => "01110111111101111100011111010001",
    708 => "01111011111111110100100110101111",
    709 => "01111001111111111100111010101011",
    710 => "01101111010101111110110010000110",
    711 => "01110110110100010110011011010111",
    712 => "01101110101110110000011100100011",
    713 => "01111111011110111000110011001101",
    714 => "01110010111011110101110111110110",
    715 => "00010111011001100111010111110100",
    716 => "01011111100111110001011000101000",
    717 => "00110010101111111000110010110010",
    718 => "01011001110111111010110011101111",
    719 => "01010111010011111111011101010110",
    720 => "01111110011111010100001000111011",
    721 => "01101011111001001100100100111001",
    722 => "01011111000101110010000011010101",
    723 => "01010101111010111100110001101110",
    724 => "01001110011011101000101001101001",
    725 => "01111111011110001110010101000100",
    726 => "01011111111101111111010101010001",
    727 => "01111111011011111111001010000011",
    728 => "01101101111101101010010000001001",
    729 => "00111110000011101100000001101011",
    730 => "01100101101101010110111001101101",
    731 => "00111011110111110101111000111010",
    732 => "00110111101101010001110101110001",
    733 => "01000110101111110110100111010001",
    734 => "01011110110100110100110100001100",
    735 => "01011111001011111110000111000011",
    736 => "01111011110111111011010111110001",
    737 => "00111101111110110110001010011111",
    738 => "01111101011111111101111010000110",
    739 => "01001000111101111001100101000110",
    740 => "01111011111111110100111100100111",
    741 => "01101010010011110111011111110101",
    742 => "01110011111101100000101101111111",
    743 => "01011101111111110110010101110000",
    744 => "01110111111101110110011011011011",
    745 => "01110111111100011101101011110111",
    746 => "01111111001111010011001111111001",
    747 => "01111111000111110000010110110101",
    748 => "00110111110011101110100100111100",
    749 => "01111101111110111001010100000011",
    750 => "01111110110111110100011010101011",
    751 => "01100111111001110110110010101111",
    752 => "01011110011111101001010111100000",
    753 => "01110011010111110100101100000101",
    754 => "00111100111110110100111101111011",
    755 => "01011010011010111000010100000000",
    756 => "01111001111001111110110111011011",
    757 => "01111111010011011110010000110110",
    758 => "01101011010110010001010110001101",
    759 => "01000111111001111111011001100001",
    760 => "01110011111011011101111011000111",
    761 => "00101111111111110101101111101011",
    762 => "00001111011111110101111000001110",
    763 => "00010101111011111111100000110111",
    764 => "01101100010110010010101011000111",
    765 => "01010011011111100011110100110000",
    766 => "01011011111101111100101111000100",
    767 => "01101111111011110100010011000100",
    768 => "01110011111110101101100011100100",
    769 => "01110011111110000111110010000011",
    770 => "01011011100101101000000001000001",
    771 => "00110001110011101100000001100011",
    772 => "01011111001101100100001111110000",
    773 => "01101110111101111010101011001100",
    774 => "01111111001111111000000000101101",
    775 => "01101111111111001001111011001110",
    776 => "01110101111011001000111101010110",
    777 => "01111001101111111110110110001010",
    778 => "01101101101111100011100101010101",
    779 => "01010100101111100000111101101010",
    780 => "01011011101111101000001110100111",
    781 => "01100100101011110111001101101110",
    782 => "01101111101110011000111100011100",
    783 => "00111110111111100010011000010101",
    784 => "01110000111101100110101100110100",
    785 => "00101101111111111100001001001010",
    786 => "01111011110111110110001001111001",
    787 => "00101111010011111011110011110110",
    788 => "00011101111111110010101000101011",
    789 => "01011101011111110001111110001101",
    790 => "00001111111111111111001110111111",
    791 => "00011010111101110000000011011110",
    792 => "01111111001110111111010110111101",
    793 => "00010101111001110100111100101111",
    794 => "00111111010111100001010001100010",
    795 => "01110110110101111101111001100001",
    796 => "01010101110111101101011101110100",
    797 => "01111101111111011011110000011100",
    798 => "01111010110011101100101101001110",
    799 => "01110111111101111000011001101010",
    800 => "01110100110010111101001110001101",
    801 => "01111011111100101010010110100101",
    802 => "01100110011000000001110111000101",
    803 => "01111101111111111001011010110100",
    804 => "00111111111110010010001100110010",
    805 => "00001110101111101011101010101101",
    806 => "00111101111011101010110011101000",
    807 => "00111101111011110001111111001111",
    808 => "01101110111100110110110100010101",
    809 => "00111111101111111001001000010011",
    810 => "01110100101111111010110110000011",
    811 => "01101111011101101100100001001011",
    812 => "00101011111011111000000011011100",
    813 => "01011111111101110010110001000011",
    814 => "01101000111111011101111111010111",
    815 => "01110101101110101010110101010111",
    816 => "01011010101111110001101111100001",
    817 => "00110100100101111000001101100100",
    818 => "01101100110011010010011000101010",
    819 => "01101110111111110001100110000100",
    820 => "01111101101110110111101101100010",
    821 => "01111010111111110000111110111111",
    822 => "01111110110011110011001101110011",
    823 => "01110101101011100010110011000000",
    824 => "01011111111100001101110000111100",
    825 => "01111011111011010110100100111101",
    826 => "01011011111111110110001110001110",
    827 => "01010110110101100000010001001110",
    828 => "01111011111111111110101010011010",
    829 => "01110011111101111100000010000111",
    830 => "01110111011110001111010001001111",
    831 => "00101110111111111100100011101010",
    832 => "00011101111111111011000111010010",
    833 => "00101101011110100010111111100011",
    834 => "01111101011111101110001001101011",
    835 => "01111110011101100001100010000001",
    836 => "00001100110101101111010110011000",
    837 => "01011110111010101101100000011100",
    838 => "01111110001010100101001011101101",
    839 => "01111011111111111100110101101110",
    840 => "00110101110111111100100101011111",
    841 => "01011111111101001000100111111001",
    842 => "01101011111111110111100011010000",
    843 => "00101110111111001101111001101110",
    844 => "00011101111111100000001110111111",
    845 => "00111011101111101001101100110010",
    846 => "01101101111010111111010110011011",
    847 => "01110101111001111100011110110011",
    848 => "01111001000111101010011111111000",
    849 => "01110000111110001110101000010110",
    850 => "01101111110101011011111101110011",
    851 => "00101011111011110111110111000010",
    852 => "01111101111111111111110111110001",
    853 => "01111011111111101100000101000100",
    854 => "01011101111011010110101101110100",
    855 => "00110101011110000101000111111010",
    856 => "01101101111111110111011001110111",
    857 => "00011011011111100001101010111011",
    858 => "00111111111101110000111000111111",
    859 => "01010011001101111010110110110110",
    860 => "01101111011111101001000011100101",
    861 => "01100111111101011000001001100010",
    862 => "01101111110111111001100111001011",
    863 => "00000101011110101101110011000011",
    864 => "01011011111001101100010000100011",
    865 => "01011111101111101011111000100000",
    866 => "00011101110001010011000010010111",
    867 => "01101110110111100101111110000001",
    868 => "01101111110110101100001001111010",
    869 => "01111101111101110110100010111101",
    870 => "00111110011110110011101101110011",
    871 => "01110111111011101101001010110010",
    872 => "01101110111111110010000100110111",
    873 => "00101111110111110001100100100001",
    874 => "01001101111110101100000010000100",
    875 => "01111100110111110001011011100100",
    876 => "01011011110111110001110100110101",
    877 => "01111011111111010010010110110000",
    878 => "01111011010110110110111000111010",
    879 => "01011011111011000101011101101110",
    880 => "01111111001011110111011010100000",
    881 => "00111111010111110100111100000100",
    882 => "01111010111101100111110110000010",
    883 => "01110111111111111000001010000010",
    884 => "01111110101111110011000110101000",
    885 => "01001101011111110001101000001010",
    886 => "00100111101110111011110111000110",
    887 => "00111011110110110110111000100111",
    888 => "01111011111110001101010111111111",
    889 => "00111001011111110111111110100000",
    890 => "01011110111001101111010100011111",
    891 => "00111111111101110101111111011100",
    892 => "01101001111111111111001011011111",
    893 => "00101101100011111101001110110110",
    894 => "01001001110100110111000110100110",
    895 => "00111110111111010100001111111110",
    896 => "01101111111101110110101110111111",
    897 => "00001011111101111100000000011010",
    898 => "00111111001111100000010011101000",
    899 => "00011011100110111111000101010100",
    900 => "01101110111110111110000100000000",
    901 => "00110111110111100000101001010100",
    902 => "01111111011101011110111010101100",
    903 => "01101101111011101100000001110111",
    904 => "00101100011101011000111001011001",
    905 => "01111011011000101011011010011010",
    906 => "01100010011111101100100000000101",
    907 => "00111101110010000111110111110010",
    908 => "01111110111111111101101110011100",
    909 => "01011111110101001110100100000111",
    910 => "01111011111101100110000010010000",
    911 => "01100001101011010100110011000000",
    912 => "01101111111111110010010101111101",
    913 => "00001101011011110101111010010000",
    914 => "01001110011110110000011101100111",
    915 => "00111011110100111100011111000100",
    916 => "01111011110011111010011011100001",
    917 => "01101111001111111110100110001001",
    918 => "00111111011111111101001111110011",
    919 => "01110111100110110011000111101111",
    920 => "00101111010110011101000010100001",
    921 => "00001001110101010010011001000011",
    922 => "01010010101111010101111000001011",
    923 => "00011100111111111110011001101101",
    924 => "01100011111011000111001000000101",
    925 => "00111011011111111100000011100110",
    926 => "01011010110111010101011010111101",
    927 => "01110101111101111010100001001101",
    928 => "01100001010111010101010001011000",
    929 => "01101111111111011000011111011101",
    930 => "00101111111011111000011110100101",
    931 => "01111101110111111011101011011010",
    932 => "01111111001011100100011010001100",
    933 => "01100110110111101100011011111110",
    934 => "01111101011011111010111101111100",
    935 => "01011111011101010111111000001001",
    936 => "01011111110110111011101110111011",
    937 => "00101101111110111000011010010010",
    938 => "01101111110111110100111101111011",
    939 => "00110101101111011011001010001010",
    940 => "01100110000011110001100101110001",
    941 => "01101111101101110011010100110101",
    942 => "01111110011111010110001010100110",
    943 => "00101001011111111111101111010111",
    944 => "01011011011101011010110010100011",
    945 => "00101110111111011100011101000111",
    946 => "00110101101010011100111010010110",
    947 => "01111101001111011010101000110101",
    948 => "01100111110111110101111010011010",
    949 => "01111001111110111111000110010111",
    950 => "00101111110111100111101001101101",
    951 => "01011101111111110111110000001101",
    952 => "01110111111011111100000111011110",
    953 => "01101111100110101000001010001011",
    954 => "01011101111100101101001101010110",
    955 => "01001011001111001001100100101111",
    956 => "01111111010011010101000011110111",
    957 => "00110110110111111011111100101000",
    958 => "00111111101111111010001001011010",
    959 => "01111111001111100111000000011000",
    960 => "01101011111010010011110001110110",
    961 => "01101101101001111100111110101101",
    962 => "01011110101110111101001110101111",
    963 => "01111110111111110011011000110110",
    964 => "01111001010111111010000100111001",
    965 => "01101111110100111101111010000000",
    966 => "01101110110110111010001110010100",
    967 => "01011111101111111010011111001100",
    968 => "01111010100101110100000100111011",
    969 => "01111101111111011101110100100000",
    970 => "01111111010111111111011101010111",
    971 => "01111011111111010100101010111100",
    972 => "00011110110000100111101101010111",
    973 => "01100011111110011001101111010000",
    974 => "01001111011111111011101101000010",
    975 => "01011101011111111110101101011101",
    976 => "01011111111110101010000000001111",
    977 => "01000111110110110001100001110101",
    978 => "01011101101100111010011110101001",
    979 => "00101111111111010110001011110000",
    980 => "00011010110100010110100000111010",
    981 => "00111101111011100100110100010101",
    982 => "01111110101011011001001001101011",
    983 => "01000011110101101010011110011001",
    984 => "01011011111100110000000101000110",
    985 => "01100011111111110000011010101111",
    986 => "00111110011010001110111011010100",
    987 => "01000111001111100001000100010010",
    988 => "01011110011111111110100001000111",
    989 => "00111111111110110010111110111101",
    990 => "01110111111111010111100101000111",
    991 => "01100111110110100100000010001111",
    992 => "00101011000101111100011010000110",
    993 => "01111111011111010110110110011110",
    994 => "01101110111101100101100111111111",
    995 => "01100001101011110111011010100000",
    996 => "01110111111101101011000110010110",
    997 => "01010111111111110001001110110001",
    998 => "00100101101001111111000001100010",
    999 => "01101110010111111110100000100111");

  constant ans_lut : lut := (
    0 => "00111000011111011101001110001110",
    1 => "01010101001010000110001000110000",
    2 => "01010100101101001101001100011101",
    3 => "00101111101100001011111011010010",
    4 => "00101111100011001110100100100010",
    5 => "00110111101101000011100100110011",
    6 => "01011010001101000110111101000100",
    7 => "01010111100111001011100100011101",
    8 => "00111010101100110111101111110101",
    9 => "01010011101101001100100010110110",
    10 => "01011010100111000001011101010001",
    11 => "00101101101010010100110101101111",
    12 => "01000111101101001101100100110000",
    13 => "01011111001010010000001000111000",
    14 => "01010110001001011100001010110111",
    15 => "01011001001011110100010000000111",
    16 => "00111001101101001110101001101010",
    17 => "01011010001000101101001110001011",
    18 => "01010100000000110111101010111010",
    19 => "00111110100011100111100000110001",
    20 => "00111110001010000110000001101001",
    21 => "01011110100110100010001000111000",
    22 => "01001001101001011111000110101110",
    23 => "01010110100110101101000001110001",
    24 => "00100110100110111001110100101101",
    25 => "01010111011111101101011101111001",
    26 => "01011011000111111011001111000010",
    27 => "00110001111101011001000000000011",
    28 => "01011110100101001110111010101000",
    29 => "00101011101101001110010101111111",
    30 => "01011011011011110010001111100000",
    31 => "01001111100110111010101001011000",
    32 => "01001111011110110100101011101111",
    33 => "00100101101101000110000001100111",
    34 => "01001100111101111100111110000000",
    35 => "01001111100101011100110001000101",
    36 => "00110001101101001011101101110011",
    37 => "01000011101100110110111000100010",
    38 => "00111010001001111000011100101100",
    39 => "00111100011111111110000100010101",
    40 => "00111000101100000001100000010110",
    41 => "00111110011110111010110000110111",
    42 => "01011010111011011001110001111011",
    43 => "00101111100011110000110001001001",
    44 => "00111100000100100101011100101000",
    45 => "01010111101011011000101100101111",
    46 => "01010010111111111010000010000100",
    47 => "01010110101101001011001110010010",
    48 => "00111111011011101110101101111001",
    49 => "01010101111011110001110000111000",
    50 => "01001101111111011000011101101000",
    51 => "01011110001100110011111011110010",
    52 => "01001100011111100010001000011011",
    53 => "00111001101101001111101011100110",
    54 => "00110111001100111101010110001100",
    55 => "00100111011110111001011001001011",
    56 => "00111101101101001110010010010001",
    57 => "00101110101100110110001011011111",
    58 => "00111010101011011101001010001010",
    59 => "00111101101100100001001100001111",
    60 => "01001111010010011100101100000100",
    61 => "00100111100111001011001100011110",
    62 => "01011110011101100010100101010000",
    63 => "01010111011110111000101010010001",
    64 => "00111111101101001010110101110111",
    65 => "00111101000111000111111101010111",
    66 => "01011011001101001101100110000100",
    67 => "01011011010111010110011011100101",
    68 => "01011100011101000110100011000110",
    69 => "01001111101011010100010100010000",
    70 => "01011110110110011110110110101011",
    71 => "01001100011011101101010011101011",
    72 => "01001110001010001011111011000111",
    73 => "01001101011111001101000010001011",
    74 => "00111110101011010100101010011010",
    75 => "00111101101100001010100111110011",
    76 => "01001111101010110111010010111000",
    77 => "01010100101101001111011110011101",
    78 => "00100011101001101111000011100011",
    79 => "01011101101101000010110111111111",
    80 => "01011110101011110000000110001101",
    81 => "01010101100111001001011010101001",
    82 => "00111110001100011111010110111000",
    83 => "01001100010001100001110110101111",
    84 => "00111101011101011001101101011111",
    85 => "01011001101001011011011010011100",
    86 => "01011110101101001000100110010111",
    87 => "00111001100110001111001000000110",
    88 => "01010110110110000101010101101000",
    89 => "01000111101101001011111111000010",
    90 => "00101111101100111101000000010010",
    91 => "01011110101010010100001111000001",
    92 => "01011100101001010101010111101110",
    93 => "00111101100011011111001100101111",
    94 => "00111010001100101101101010101100",
    95 => "01001011101100110101011001100011",
    96 => "01000010010111001010000011111101",
    97 => "01010110001011000001101001000101",
    98 => "01001011100110010001010010001110",
    99 => "01011011101100100010000110000011",
    100 => "00101101100100010110110011011111",
    101 => "00101110101010010010110001101011",
    102 => "00111111100110100110000111111100",
    103 => "01001100100111000001100001100101",
    104 => "01010000101100100111111110110100",
    105 => "00110010001100011101101110100001",
    106 => "00101111100001110111011010100111",
    107 => "00101111100111001010000110110100",
    108 => "01001001101100001011001101000011",
    109 => "00111111011100101001010111010001",
    110 => "01001110101101001111101011101110",
    111 => "01011011101000000111000001010100",
    112 => "01011110101100011101110110110011",
    113 => "01011101100110101110010100011111",
    114 => "01011011100111111010111101110101",
    115 => "01011110101101000100010001110010",
    116 => "01011011001010010101011000100111",
    117 => "00111101011111111111010100110101",
    118 => "01010101101011100111100010010010",
    119 => "01011111011011101011110110100001",
    120 => "00111111011111111111011000111011",
    121 => "00111100101101001011101000000110",
    122 => "00100111101011101000100011011101",
    123 => "01001111101100100000101001111000",
    124 => "01011011011110011011010111010000",
    125 => "01011101100001111010000111011001",
    126 => "01011111000111000111101000011000",
    127 => "00111110011001110000001000101111",
    128 => "01010101000101111000101011110111",
    129 => "01011011011111111110101111001001",
    130 => "01001100110111110001111111110010",
    131 => "01011110001011011011100011011010",
    132 => "01011010001001111001000111011001",
    133 => "00110100001011110000010001010101",
    134 => "01011110101101001010111001010011",
    135 => "01011011100011100111100010001001",
    136 => "01011111001101001100111010000111",
    137 => "00111101100110010100011111001100",
    138 => "01011011000111110100010011011111",
    139 => "01001111101010001111010100101000",
    140 => "01011011101101000010011010000111",
    141 => "01010111101100110111101110010001",
    142 => "00101011011011010011010011111111",
    143 => "01010110101011111101101001111001",
    144 => "00110010101100001111110100101100",
    145 => "01000011100111000101111011001110",
    146 => "00111100001010011101011111100010",
    147 => "00100101101010001010000111110100",
    148 => "01011101101010011011111100100010",
    149 => "01011111001011101110100101000010",
    150 => "00101011101101001011101001001101",
    151 => "00110110011111111111100100100001",
    152 => "01010111101001110010111000100110",
    153 => "01011111011111101111100100101001",
    154 => "01001110100011101111101111011001",
    155 => "00111111101101001110101001000110",
    156 => "01001111100110111011000111101010",
    157 => "01010111101100100001010101001100",
    158 => "00101101001011011111111110000010",
    159 => "01001010101010000100000101110000",
    160 => "01011101101101001110101001101001",
    161 => "01010111001001110110110111101110",
    162 => "01011111011111111101001101100001",
    163 => "01001111100110010101001001110110",
    164 => "01011111001100011110001000001011",
    165 => "01011011100011101101101001101101",
    166 => "01010111011010010001010011111010",
    167 => "01010110111101011000011111001010",
    168 => "00111111101101001100110110111011",
    169 => "01011011101101000101110011100101",
    170 => "01010111001100110000010110011110",
    171 => "01011111010111010011011110110110",
    172 => "01010110011011100000011111000010",
    173 => "01001010100011011100011010011011",
    174 => "01011011001010010100110010001000",
    175 => "00110001101100110000001000110001",
    176 => "01011111000111001000011111000101",
    177 => "00111101101101010000001010010111",
    178 => "00110111010111010011100000110011",
    179 => "01011110011110101000011010011011",
    180 => "00110110101100110101000001000111",
    181 => "01001101100110111001001110111111",
    182 => "00110110101100100000000011110111",
    183 => "01010111000111000011011011001010",
    184 => "01010011011111111101010000011010",
    185 => "01010111001010010010110000011000",
    186 => "01010110010010111000101101110000",
    187 => "01011110000111001010000101110010",
    188 => "01011110101100111100001001011110",
    189 => "00111111001100111110000010001110",
    190 => "00101111101101001010001100101111",
    191 => "00110111101101001111000110101101",
    192 => "01011101101101000101010111001111",
    193 => "00111101010110010000010101100110",
    194 => "00101111001011001110011110101000",
    195 => "01011011101010010100000000001010",
    196 => "01001111011110011011110001000111",
    197 => "01011011001001010100110001110111",
    198 => "01000011001100011111011110111100",
    199 => "00111111001100100111111000001001",
    200 => "00111101001101000100101011100100",
    201 => "00111111100101011010110011110010",
    202 => "01001010001111110110000010010010",
    203 => "01010110000110111011001011110011",
    204 => "01001100101010000011101110010101",
    205 => "01010100101101001011001101111111",
    206 => "00110101001010010011110111110001",
    207 => "01010100111101110100001000010011",
    208 => "01010100101100011111110000011010",
    209 => "01011101101100111001111010010111",
    210 => "00101111101001100011001111111101",
    211 => "01011011011011110001100110111001",
    212 => "01001110011101011001001111010100",
    213 => "01011101000111001000111011001111",
    214 => "01001011001011011000001010110011",
    215 => "00110111101011100010100111110100",
    216 => "01011111001001111011100101111010",
    217 => "00100111101101010000010001111111",
    218 => "01000111010111001001101000011001",
    219 => "00111101011101111011011000000100",
    220 => "01001111101100010100001111100011",
    221 => "01011101101010001111001111001001",
    222 => "00110111011100110000010110100010",
    223 => "00111110000111000101110111011101",
    224 => "01010111101101000101111100010011",
    225 => "00111011001100001011011100110111",
    226 => "01011110101101001011000000010100",
    227 => "01011111010011100111111101000111",
    228 => "00110111001101001101101000010010",
    229 => "00101111101001100010010010100000",
    230 => "01010011101011101101110001110000",
    231 => "01000111011111111101001100010100",
    232 => "00111111000000110001100000001110",
    233 => "01011111001011010111001011100011",
    234 => "01010101001100010111100000001011",
    235 => "00111110011001000100111100001100",
    236 => "01000110101100000101111111101001",
    237 => "01010101101011001010000111111001",
    238 => "00101011101010010100000010001001",
    239 => "01011010111111011101111011111111",
    240 => "01011101100110100000011111111110",
    241 => "00111010011101111001010000100110",
    242 => "01011110100101011110010011101110",
    243 => "01001111001100001001011000011011",
    244 => "00101110101100110111110011111011",
    245 => "01001110001100100000111110111100",
    246 => "00100111011111011010100010010100",
    247 => "01010111101100011101000101110001",
    248 => "01001101101001111111101111001100",
    249 => "00111110110001001011011001000010",
    250 => "01011100010010010000000000000010",
    251 => "00101111101100011110100110110100",
    252 => "00111101101100111000010000001011",
    253 => "01010111010101011100011000101111",
    254 => "01011110100110111101101100000010",
    255 => "01010111101101001010011111101110",
    256 => "01001011001100001000000000101011",
    257 => "01011110101100100001101001110000",
    258 => "00111111011010101010010100110100",
    259 => "01011001101011110000001111001101",
    260 => "01011100111110101100110100111001",
    261 => "00111111011011110010100110000010",
    262 => "01000011101101001011101000110000",
    263 => "00101100100101111001011111011010",
    264 => "00111111000110100010111001000001",
    265 => "01010010011111110001110011110110",
    266 => "01011111011111010100111010001000",
    267 => "01001110101100110100110110101111",
    268 => "01011100111010110111000101010010",
    269 => "01001100011011000101010000011011",
    270 => "00100011011011001101111010001000",
    271 => "01010111101100110101010100101010",
    272 => "00111111101101001101111010101100",
    273 => "00110111101011101001111010010101",
    274 => "00111101101101010000010001101000",
    275 => "01011111001000001011000011000010",
    276 => "01010110101001111100110111100111",
    277 => "00110111101100111000010001111000",
    278 => "01011010101100110100101011010001",
    279 => "01011110111010100111111010110100",
    280 => "01011101101101001010110001011100",
    281 => "01001001011011110101001110000001",
    282 => "01011110101001000011101001111101",
    283 => "00111111010011110001000000100100",
    284 => "00111011011111111011000011011011",
    285 => "01011010101101010000001000101010",
    286 => "00110111101101001010000100001111",
    287 => "00111110010010110000110010110001",
    288 => "01011101101101001110111111101111",
    289 => "01010110101100101011110111011011",
    290 => "01011010111111111010001111011111",
    291 => "01001111100101010000001101001100",
    292 => "00111111101101001010110101110010",
    293 => "01001101100111001011010010011010",
    294 => "01001111011110111111010001111011",
    295 => "01001101010100100010011101110101",
    296 => "01011101101011111101011110100111",
    297 => "01000011101011001111000010011111",
    298 => "01011110011111111101100010000010",
    299 => "01000111100101010011110000011101",
    300 => "00111111001000110000001110000101",
    301 => "00110111101001010100111001101010",
    302 => "01011011000111001100000100110110",
    303 => "01001011101100010010010000000100",
    304 => "01011111001100110111001001010111",
    305 => "01011101100110100000000001011010",
    306 => "01001111101011101001101011000001",
    307 => "01011110000110100110110010011110",
    308 => "01001010101010010101000011111000",
    309 => "01011101100101101000111010111010",
    310 => "00111110001011110011101100110111",
    311 => "01011011101010010100001000011100",
    312 => "01011111000111000110101100110001",
    313 => "01010110111111111101001001111100",
    314 => "01011100111111110101101001111101",
    315 => "01011101011111111100110101110010",
    316 => "01001101011100110101010000110001",
    317 => "01011001101001111010000000000011",
    318 => "01010101101100111000100111001111",
    319 => "00111100101100011111111001011101",
    320 => "01010000001101000000100011010110",
    321 => "00100110101010101001010001010110",
    322 => "00111011111011010000001011101100",
    323 => "00100101101001111001111101000110",
    324 => "00111111101101001010111001010011",
    325 => "01011011010111010111101001000000",
    326 => "01010001100011101110010111111001",
    327 => "01011101101101001000111110000011",
    328 => "01011001010100111111101111000000",
    329 => "00111001101011101110100000010110",
    330 => "01010110100001111010111111110010",
    331 => "01011100100110110111010100100011",
    332 => "01010110101011101100001010110011",
    333 => "01010111100011101011100110001110",
    334 => "01011111011111111001011010011000",
    335 => "01010111101100010111001101010001",
    336 => "01011011100111000111010111111010",
    337 => "01010111011011110000001000001111",
    338 => "01011011101010000110011000101011",
    339 => "00101110101001101010110011001111",
    340 => "01001111100010110100101111010110",
    341 => "01011110101010010100110111010110",
    342 => "01001100101011010101111000100001",
    343 => "01010111011100100111000111101001",
    344 => "00100101100100011111100101111000",
    345 => "01010110101100110000100011001101",
    346 => "00111111100111001000111110000101",
    347 => "01011101101101001011001011011000",
    348 => "01011100010010100001001110110000",
    349 => "01011110001101001011000001010111",
    350 => "01011110101101000010101001100111",
    351 => "00111101101011001011110000001011",
    352 => "01011010011111011011110010110110",
    353 => "01001110101100110111001011101001",
    354 => "01011010111111011011000101110010",
    355 => "01011111011111100110010100101010",
    356 => "01011111001101001011101001100010",
    357 => "01001100101001110010111010000010",
    358 => "01010101111111111000000011011110",
    359 => "01001101001001101111011110100011",
    360 => "01011110100011110000000001001110",
    361 => "01001011001101001101111000100100",
    362 => "01001011100101011101111010011010",
    363 => "01011110101100101111010100000101",
    364 => "01011011101001011110000001110001",
    365 => "01001100101100001101000100001101",
    366 => "01001111010100111010011010101111",
    367 => "01011101101100110100110101100101",
    368 => "01001111101101001011001100011110",
    369 => "01010110101100110111100000000000",
    370 => "01011101011001100011000010001011",
    371 => "01010001001101001111100101101101",
    372 => "01011011101101001010100011100001",
    373 => "00110110001100111000011100111100",
    374 => "00111101101100011000100101110101",
    375 => "00100100101100010110111001011100",
    376 => "00101111011111110101110001111101",
    377 => "01001101101100110110000000000010",
    378 => "01000110010010011111101001110100",
    379 => "01001101010100111000001111101001",
    380 => "00111111101101000001010101100001",
    381 => "00111011101100110110011011111110",
    382 => "01010111011111011011100101001011",
    383 => "01010111101100010111011011000000",
    384 => "01011001001101001101100101100000",
    385 => "01011110101001000110100000011001",
    386 => "01011111001011101100000001101000",
    387 => "01011101110001111000111011110100",
    388 => "01011011001100011000111010110000",
    389 => "00100101100101001111110111100110",
    390 => "01011110101011100101110111010101",
    391 => "01011111000110011010110100000110",
    392 => "00101111001000100111110000001011",
    393 => "01010110100111001011101000011111",
    394 => "01011011011111111000001001111001",
    395 => "00100111101011110011000100001000",
    396 => "01001011011110111001000010010110",
    397 => "01010111101100101011010110011001",
    398 => "01010011101010111110011000011010",
    399 => "01011100101001111001010010001010",
    400 => "01011101101001011111111111011000",
    401 => "01011111010110110101100000001110",
    402 => "00110111101000110010101001101111",
    403 => "00110011001000010111001100001000",
    404 => "00110111101101001110010010011100",
    405 => "01011111001100010101110011010111",
    406 => "01001010001011101110100111010110",
    407 => "00101011101011101011001011000011",
    408 => "00111011001101001110000101110101",
    409 => "00111111101100001010010001111100",
    410 => "01010111101101001100010011110100",
    411 => "01001100001101001011110011000000",
    412 => "00110111000100111100111110011000",
    413 => "01011101101000100110011101000100",
    414 => "01010111100110111001001101010111",
    415 => "01011100001101001101101100111001",
    416 => "00110010101100101110010001101011",
    417 => "01001110001000100010010111010001",
    418 => "01011100100000111100000001100010",
    419 => "01011011011000011110010010000110",
    420 => "01010101101100011100011010101110",
    421 => "01001001101101001101000111001111",
    422 => "00110111101101000100000100101110",
    423 => "01010010101101001110001001011101",
    424 => "01010001001101001101101000110111",
    425 => "01001011101001110101000101111001",
    426 => "01001111100110101001101011100101",
    427 => "01011101101010001100101001111011",
    428 => "01011111010001110110000010111001",
    429 => "01011001101010010010010110011000",
    430 => "01010110110111010011100000000100",
    431 => "01011101100110100111001010111111",
    432 => "01011101101101000101111110000000",
    433 => "01000110100111001000010100001010",
    434 => "01011011101011100010000101100111",
    435 => "00111111001101001101000111000000",
    436 => "00111011101101000111000001100100",
    437 => "00111011101100110110100111101000",
    438 => "01011010100110100111000100111010",
    439 => "01011110101101000011000000110111",
    440 => "01010110101100011111011101100101",
    441 => "00111011101101001101100100111100",
    442 => "01010011101100001111011101100010",
    443 => "01011110101100011001100011111001",
    444 => "01010001101000010101110100001101",
    445 => "01011011011011110100110100101110",
    446 => "01011111011110110111101011010001",
    447 => "01011011101010000101111110111111",
    448 => "00110101111110111000111101111100",
    449 => "01011101011111011000000011000110",
    450 => "00111111101011100011000100110101",
    451 => "00110110111011100101111100011101",
    452 => "00111111101100010101111011010110",
    453 => "01001101111111011011101100010111",
    454 => "00101111001001111111110011100011",
    455 => "00111111101100111111100001001110",
    456 => "01001111001011100100100101111010",
    457 => "01011101101010111111101101011101",
    458 => "01011001011111111101011111100000",
    459 => "01011100111100110011100001101010",
    460 => "01011111011001010110011000100100",
    461 => "01011011010110000010110000101011",
    462 => "01011110101010010100110100100100",
    463 => "01011000101000110001001010110010",
    464 => "01011111011110111010101100110111",
    465 => "01000011101011010111101100111111",
    466 => "01011100111101000101101011111000",
    467 => "01001111101100010011101010010111",
    468 => "01010100100111000110110000110100",
    469 => "01010111101101001101110001010110",
    470 => "01011101100011010001111100111001",
    471 => "01011100111111111011100010010001",
    472 => "00101011011111001101000011111101",
    473 => "00111110101001010011000000101010",
    474 => "01011111001101001011011011001110",
    475 => "01010010100110111000110111111000",
    476 => "01010011101101000000011100101111",
    477 => "01011101100011011100111101111001",
    478 => "00100101101011110011100001111110",
    479 => "01011101100101011100100101011110",
    480 => "01011110001100010011101110101101",
    481 => "01011001011111110101000101100100",
    482 => "01010111011110001000111101101100",
    483 => "01001111001101001111100010011001",
    484 => "00101110100110111111100111100010",
    485 => "00110011001101001100101001011011",
    486 => "01011001011010111000110011101111",
    487 => "01000111101101001100000001010110",
    488 => "00111110111111111011000110101010",
    489 => "01011101101001110100000001001101",
    490 => "01011111001101001011100110010010",
    491 => "01011011100010010110101111100010",
    492 => "01011011101101001101010100011100",
    493 => "01011111010101111111111100100100",
    494 => "01011111000111001000011000101110",
    495 => "00110100101100110100000111010011",
    496 => "01001100001101000101100010110101",
    497 => "00111101101001011111100000001101",
    498 => "00111101111111111010110100000100",
    499 => "00101101100110111110000011111000",
    500 => "01001110101100110100100110111101",
    501 => "01000111101010010010001001010010",
    502 => "01011111000111001001000001011101",
    503 => "00101011100110010011000010111000",
    504 => "00111101011011001101100110110110",
    505 => "00101111100110010101001010000100",
    506 => "01011101100101100000010101100000",
    507 => "00110111101011111010010010000110",
    508 => "00111110011110111100110110110111",
    509 => "01011111011000100001101101010100",
    510 => "01011011001011111010011010111010",
    511 => "01000001001001110111011001111000",
    512 => "01011111001011101001111100101000",
    513 => "00101111010111001111000100011101",
    514 => "00101101011001010011011011010000",
    515 => "00111111101001100011101110101001",
    516 => "01010111100101011110110110100010",
    517 => "01011010001100111010111110000001",
    518 => "01001101011101110110010101010100",
    519 => "01001111101011110010110011110110",
    520 => "01011111000001110110100110100011",
    521 => "00111101101001100000001000100111",
    522 => "00111101011110110111100001011001",
    523 => "01011111001000110010001010110101",
    524 => "00111010101011110011010110000111",
    525 => "01010111101101001010011111010011",
    526 => "01011111001101000100100001010110",
    527 => "00110111011111101111111011101111",
    528 => "00101001101001100010001100000101",
    529 => "01011110101001011111010110010011",
    530 => "01011110100110110000000110001101",
    531 => "01011101101101000000010101110100",
    532 => "01010001101011111100010110110000",
    533 => "01011100101010010010010100001110",
    534 => "00111111101100011100111101011100",
    535 => "01011001101000010011111100000111",
    536 => "01010101011101010110001000110010",
    537 => "01010001001001000000000101010111",
    538 => "00111111011101010011010000000111",
    539 => "01010010101101001110000111110000",
    540 => "00111110110111000110111110110011",
    541 => "01000111001011011000110001000111",
    542 => "01011110011000101101110011011110",
    543 => "01011110011100000000011011010010",
    544 => "01011111011111110111011100001110",
    545 => "00101111101101001010110110101010",
    546 => "01010111101011011011111100010000",
    547 => "01010000011010010111111011000100",
    548 => "01001110101100111111100100010111",
    549 => "00111011011111111011010111100100",
    550 => "01011101101101001101000101010100",
    551 => "01011101111111100010000010010101",
    552 => "01001101101000101100111111101000",
    553 => "01001010101100111011111111101100",
    554 => "00111011011010100000101111110111",
    555 => "00111011011111111111101001101111",
    556 => "01010001101101001100111110010011",
    557 => "01011111001011110011011101010110",
    558 => "01010110110111011010111000010010",
    559 => "00100111100110100101010111010010",
    560 => "01010101101100111000111001111011",
    561 => "01011011100111001011000110111101",
    562 => "00110101100110101010001110100000",
    563 => "00111111100011010000000001010100",
    564 => "01010111101101000111000101011100",
    565 => "01011110101100011111101110111111",
    566 => "00111111100011101100111111001001",
    567 => "01010001101101000110001110010011",
    568 => "01011011101100101111001011011101",
    569 => "01011111001100011111111010011100",
    570 => "01011100101001011101110001010001",
    571 => "00101101000101000000001101000101",
    572 => "01010011101010010001100011000010",
    573 => "01011110010010100000101101100000",
    574 => "01000111100010100010011010100101",
    575 => "01001110100100100010010101101011",
    576 => "01010101100011101111011110101100",
    577 => "00101111101100110101110100111101",
    578 => "01010011000101000111010111100011",
    579 => "01011011101101000110101110101101",
    580 => "01001010001000100101010010111001",
    581 => "00111001011011100000101001101000",
    582 => "01011101101100010001111010010100",
    583 => "00101011011011101111010010100111",
    584 => "01001111011011000110001111111010",
    585 => "00110011101011100001100110000000",
    586 => "01011111001011011010010010010111",
    587 => "00110101111101110111001101001110",
    588 => "01010111001011000000001100011011",
    589 => "01010011101100110100100110111101",
    590 => "01011011100011101110000110001000",
    591 => "00101111100001111110011011000010",
    592 => "01001110011001010100010110100100",
    593 => "01010111001100110010101100101011",
    594 => "00101110011110111111000010000010",
    595 => "00101101101010010011010110010000",
    596 => "01011100101011011111001010100001",
    597 => "01011111001000010100011001001010",
    598 => "01011111001000011111100110110011",
    599 => "01010010101011110011100101110001",
    600 => "01011110011111110000110100001011",
    601 => "01010010100111001010110000101111",
    602 => "01011101011111101000110000010001",
    603 => "01010110100000110001011000101111",
    604 => "01001111011111110010001001001101",
    605 => "01010011101000101011111111010101",
    606 => "00111110101011110000011001111101",
    607 => "01011111000110101101111000110110",
    608 => "01011011100100101110001000100101",
    609 => "00111101100111000010100011010101",
    610 => "01010101011110101100110001101010",
    611 => "01011011101101001010101100101111",
    612 => "01001011101010010000111010101110",
    613 => "01010110001100100001011001110110",
    614 => "00110011000111000000110011101111",
    615 => "01011110101011110010110100110011",
    616 => "00101101001100101111100111111111",
    617 => "01001111100101101110101101101100",
    618 => "01011110100110001001010111101101",
    619 => "01011001001011000001110011001101",
    620 => "00101101001101001111110010011100",
    621 => "00110101101101001011100111001010",
    622 => "01001111101100110100111111010100",
    623 => "01011011100001101011111000000111",
    624 => "00111101001011110011001100001100",
    625 => "01001111101011110000111110010010",
    626 => "00100100101011110011001011000010",
    627 => "01011011001010010010100100001111",
    628 => "01011001100110000010100011000010",
    629 => "00111111101100110101000110000111",
    630 => "01011111000111000001001010001111",
    631 => "00111110011111011011010100110100",
    632 => "01011111001100111101101011010010",
    633 => "00111101101011011000101000011010",
    634 => "01011111001001000100001010111111",
    635 => "01000110101011110010010011101110",
    636 => "01010100111011101111101010000010",
    637 => "01000001001101001011110100110111",
    638 => "01011101001101001011111010010101",
    639 => "00101110111110110001000000010110",
    640 => "01011111010111011010111001000110",
    641 => "01011001001101001010010101000000",
    642 => "01011011101011110000001101001010",
    643 => "01011010101011001101100100101110",
    644 => "01011101011111111000011111101010",
    645 => "01011110011001111111101000111000",
    646 => "01001001000110110000010001011110",
    647 => "00101111101010000110000111110110",
    648 => "00101110101101001101111000111011",
    649 => "01010011101010010000000111010101",
    650 => "00111011101100100000001000100101",
    651 => "01010010000111001000111010011011",
    652 => "00111111010011000110010110100100",
    653 => "01010011001100110100000110101110",
    654 => "00111101101100010111010111011000",
    655 => "01011101001001010111101101010100",
    656 => "01001111001101001101001011101101",
    657 => "01011010101101100011001100010101",
    658 => "01011010101001100011010000000011",
    659 => "01011110001101001110100011111101",
    660 => "01000101101100111001010111110000",
    661 => "01001110101101001111000011000101",
    662 => "00110110111111011001011101101001",
    663 => "00111111001011110100010010010010",
    664 => "01000011011001000000111000110100",
    665 => "00101111011111011110100010100101",
    666 => "00111111000100110001011001001111",
    667 => "01001111011100110100110111000000",
    668 => "00111001100100001101010001111010",
    669 => "01010001101010000111111000001101",
    670 => "00110100100001010010100011101000",
    671 => "01011110101010101000011010011111",
    672 => "00100001100111001001101011100111",
    673 => "01011110100110111000001001011001",
    674 => "01011010100110001110111100100110",
    675 => "00111111011000001101110111101010",
    676 => "01011111000110101110000001111100",
    677 => "00111001110010011101000100011000",
    678 => "01010111100101011110010110111110",
    679 => "00110111101101001100010011110101",
    680 => "00111101101010000101111111100011",
    681 => "00111111100111001010000010000110",
    682 => "01011111011111011101101100011100",
    683 => "01011111011001101000001100001100",
    684 => "01011111001011101011101110001011",
    685 => "01011111011110101010010100100010",
    686 => "00111110101010101001010100110010",
    687 => "01001011101101001111101100011000",
    688 => "01001111101101001011000000110010",
    689 => "01000111100011011110010100010000",
    690 => "01011111010110001101111001001000",
    691 => "01010111100111000101010010110101",
    692 => "01011100101100110110100100101000",
    693 => "00111101010001010100101011101000",
    694 => "01001111100011101100110100111110",
    695 => "01011011011111000100001011101010",
    696 => "01011010011111011000110110110011",
    697 => "01000110100111001000100101001110",
    698 => "01001110101001111010000100000110",
    699 => "00111111100100111111110110111100",
    700 => "01000111101011011001100111100101",
    701 => "00101101100001111010011101011100",
    702 => "01000101001100110111010011111110",
    703 => "00110111011011101101111001101100",
    704 => "01011101101101001110100100101001",
    705 => "00111110011101111000111101101101",
    706 => "01011101101100010011110100101001",
    707 => "01011011101100100001011011101111",
    708 => "01011101101101001100010001110010",
    709 => "01011100101101001111001110000001",
    710 => "01010111011010110001110000001110",
    711 => "01011011001000111011011110101101",
    712 => "01010111000110101011100101100011",
    713 => "01011111011111011100001111100111",
    714 => "01011001001011110000101000111000",
    715 => "00101011011100101110010100011010",
    716 => "01001111100011101011001100000010",
    717 => "00111001000111001001010101010110",
    718 => "01001100101010010011010010010100",
    719 => "01001011011001101011110010001011",
    720 => "01011110111111101010000000101011",
    721 => "01010101101010110010000010100001",
    722 => "01001111010001001011000111011011",
    723 => "01001010101011011011101011110100",
    724 => "01000110111101110001110110111110",
    725 => "01011111011111000110110000111011",
    726 => "01001111101100100010011101001001",
    727 => "01011111011101111101011111111101",
    728 => "01010110101100011010110111110101",
    729 => "00111110101111110010101001111100",
    730 => "01010010100110000110010001000010",
    731 => "00111101101010010001011011001100",
    732 => "00111011100110000100001000111011",
    733 => "01000011000111001000011100010100",
    734 => "01001111001001000111010101010000",
    735 => "01001111010101000011000101010111",
    736 => "01011101101010010011011111111101",
    737 => "00111110101100110110000101011110",
    738 => "01011110011111111110111101000010",
    739 => "01000100001100100000011000110101",
    740 => "01011101101101001100011001100001",
    741 => "01010100111001100111010111010111",
    742 => "01011001101100010111011011111011",
    743 => "01001110101101001100111001000101",
    744 => "01011011101100011111010000010100",
    745 => "01011011101011111111001010000111",
    746 => "01011111010111000001010011101100",
    747 => "01011111010010011100010000110111",
    748 => "00111011101000101011110110101110",
    749 => "01011110101100110111001101010111",
    750 => "01011111001010010000110111100010",
    751 => "01010011101011000001110010000110",
    752 => "01001110111111110100101010101111",
    753 => "01011001011011110001011001111111",
    754 => "00111110001100110101101010001001",
    755 => "01001100111101011000101111011100",
    756 => "01011100101011000100110010000111",
    757 => "01011111011001011001010100101010",
    758 => "01010101011010111011110110001100",
    759 => "01000011101011000100111110110010",
    760 => "01011001101011100111110111100110",
    761 => "00110111101101001100101011100110",
    762 => "00100111011111111010111011111001",
    763 => "00101010101011110100001010010110",
    764 => "01010101111010111100100100010010",
    765 => "01001001011111110001111000110100",
    766 => "01001101101100100001100001011011",
    767 => "01010111101011110000000100000010",
    768 => "01011001101100110011000000110011",
    769 => "01011001101100100101011111010100",
    770 => "01001101100010101100101110010110",
    771 => "00111000101000101010110110011101",
    772 => "01001111010110000000001001010101",
    773 => "01010111001100100000110010000010",
    774 => "01011111010111010110100111111111",
    775 => "01010111101100111101001000001010",
    776 => "01011010101011100000001010110010",
    777 => "01011100100111001011110011100110",
    778 => "01010110100111000000101001100100",
    779 => "01001010000110111111100100110001",
    780 => "01001101100111000010100011011100",
    781 => "01010010000101011101101111100101",
    782 => "01010111100110100001110110001010",
    783 => "00111111001101000101110100010110",
    784 => "01011000001100011001100101111011",
    785 => "00110110101101001110111100100000",
    786 => "01011101101010010001100001101000",
    787 => "00110111011001101001110000100111",
    788 => "00101110101101001011100101001001",
    789 => "01001110011111111000111110101101",
    790 => "00100111101101010000000010011101",
    791 => "00101101001100011100111101100010",
    792 => "01011111010110110101101110001001",
    793 => "00101010101011000001000110001101",
    794 => "00111111011011100110111111110111",
    795 => "01011011001001100011100111101111",
    796 => "01001010101010001110001111000010",
    797 => "01011110101101000011011101111000",
    798 => "01011101001000101011000111101001",
    799 => "01011011101100011111111101101101",
    800 => "01011010001000011000010111110110",
    801 => "01011101101100000011110000110001",
    802 => "01010010111011111000011100111000",
    803 => "01011110101101001101111110110100",
    804 => "00111111101100101001001110011010",
    805 => "00100111000111000011111101101000",
    806 => "00111110101011101100100101110000",
    807 => "00111110101011101111001101111110",
    808 => "01010111001100001000010010001111",
    809 => "00111111100111001001011110001001",
    810 => "01011010000111001010001010111111",
    811 => "01010111011110110101100101010100",
    812 => "00110101101011110001011011111011",
    813 => "01001111101100011101111100000000",
    814 => "01010100001101000100010000101000",
    815 => "01011010100110101001010000111001",
    816 => "01001101000111000110011100110011",
    817 => "00111010000010110100001011100000",
    818 => "01010110001000100000101111101001",
    819 => "01010111001101001011001101100011",
    820 => "01011110100110101110100101110001",
    821 => "01011101001101001010111111101101",
    822 => "01011111001000101101101011011011",
    823 => "01011010100101010101000000100000",
    824 => "01001111101011111001010111000110",
    825 => "01011101101011100101001011000100",
    826 => "01001101101101001100110110011010",
    827 => "01001011001001011000001100000100",
    828 => "01011101101101001111110101100001",
    829 => "01011001101100100001010001010001",
    830 => "01011011011111000111001111011100",
    831 => "00110111001101001111000101111000",
    832 => "00101110101101001110100101001100",
    833 => "00110110011111010001001110101011",
    834 => "01011110011111110111000100001101",
    835 => "01011110111110101111111110111110",
    836 => "00100110001001011110000000110111",
    837 => "01001111001011010110000011011011",
    838 => "01011110110100001101000000101001",
    839 => "01011101101101001111001100010000",
    840 => "00111010101010010011111101010110",
    841 => "01001111101100001110101110111100",
    842 => "01010101101101001101010100100000",
    843 => "00110111001100111110100010101101",
    844 => "00101110101101000101000011100111",
    845 => "00111101100111000011001010000010",
    846 => "01010110101011011100101000011110",
    847 => "01011010101011000011111001011010",
    848 => "01011100010010011000100010110101",
    849 => "01011000001100100111111100100001",
    850 => "01010111101001010110100001100010",
    851 => "00110101101011110001010111011001",
    852 => "01011110101101010000010000111000",
    853 => "01011101101101001001010000011111",
    854 => "01001110101011100101001110010100",
    855 => "00111010011111000010000110000000",
    856 => "01010110101101001101010001001100",
    857 => "00101101011111110000110011101001",
    858 => "00111111101100011101010000110011",
    859 => "01001001010110001101100001001011",
    860 => "01010111011111110100100000110000",
    861 => "01010011101100010100010110000010",
    862 => "01010111101010010010110101010111",
    863 => "00100010011111010110101100001011",
    864 => "01001101101010111101110111001110",
    865 => "01001111100111000100000011010001",
    866 => "00101110100111101101111100110111",
    867 => "01010111001010001011011001000111",
    868 => "01010111101001110101010111110000",
    869 => "01011110101100011111010011000001",
    870 => "00111110111111011001101011011011",
    871 => "01011011101011101101011101000110",
    872 => "01010111001101001011011000011101",
    873 => "00110111101010001111110010100011",
    874 => "01000110101100110010011101111111",
    875 => "01011110001010001111101111001010",
    876 => "01001101101010001111111000101110",
    877 => "01011101101101000000001000000101",
    878 => "01011101011011010000001011010010",
    879 => "01001101101011011110111000100001",
    880 => "01011111010100111111000010101100",
    881 => "00111111011011110001100010100011",
    882 => "01011101001100011010000000010100",
    883 => "01011011101101001101100010001111",
    884 => "01011111000111000111000000011100",
    885 => "01000110011111111000110011101010",
    886 => "00110011100110110000010011011100",
    887 => "00111101101001111001011110001100",
    888 => "01011101101100100111011111101101",
    889 => "00111100011111111011111111001000",
    890 => "01001111001010111111000000001010",
    891 => "00111111101100011111000110010000",
    892 => "01010100101101010000000001001110",
    893 => "00110110100001111010111011010011",
    894 => "01000100101001001000001110001110",
    895 => "00111111001101000000110011001011",
    896 => "01010111101100011111010111010110",
    897 => "00100101101100100001010000101010",
    898 => "00111111010111001000111001001111",
    899 => "00101101100011010100100000111111",
    900 => "01010111001100111000111001101111",
    901 => "00111011101010001001010111110101",
    902 => "01011111011110101110101001101000",
    903 => "01010110101011101101000010011010",
    904 => "00110101111110101011100101000000",
    905 => "01011101011100001110100101111010",
    906 => "01010000111111110110001111010010",
    907 => "00111110101000000011001001011000",
    908 => "01011111001101001111100000010100",
    909 => "01001111101001010001010101010110",
    910 => "01011101101100011001010110100110",
    911 => "01010000100101001110111111111110",
    912 => "01010111101101001011011110100000",
    913 => "00100110011101111000101110001001",
    914 => "01000110111111011000000010010100",
    915 => "00111101101001001010010100001011",
    916 => "01011101101000110000100000110010",
    917 => "01010111010111011010011011011110",
    918 => "00111111011111111110100111111000",
    919 => "01011011100011001111000101110000",
    920 => "00110111011011000010001100001010",
    921 => "00100100101001010010110100010001",
    922 => "01001001000110111011000001011000",
    923 => "00101110001101001111101111100111",
    924 => "01010001101011011111011111101001",
    925 => "00111101011111111110000001110001",
    926 => "01001101001010000101000110111001",
    927 => "01011010101100100000101110011100",
    928 => "01010000011011100000100011001001",
    929 => "01010111101101000010010011101001",
    930 => "00110111101011110001100101110110",
    931 => "01011110101010010011100111011000",
    932 => "01011111010100110011100010110111",
    933 => "01010011001010001101110110000101",
    934 => "01011110011101111011010101011101",
    935 => "01001111011110101011000011101101",
    936 => "01001111101001111011010100101010",
    937 => "00110110101100110110111000110001",
    938 => "01010111101010010001000100110111",
    939 => "00111010100110111101001100010001",
    940 => "01010010101111110110011000001101",
    941 => "01010111100110010010001011001010",
    942 => "01011110111111101011000001110110",
    943 => "00110100011111111111110111101011",
    944 => "01001101011110101100100010110110",
    945 => "00110111001101000011101101101111",
    946 => "00111010100100110110110111001110",
    947 => "01011110010111000101100110100101",
    948 => "01010011101010010001011011110001",
    949 => "01011100101100111001010001011001",
    950 => "00110111101010001100000001111110",
    951 => "01001110101101001101011001000110",
    952 => "01011011101011110010111010111101",
    953 => "01010111100011001010000110110110",
    954 => "01001110101100000100110011001000",
    955 => "01000101010110111011101011010011",
    956 => "01011111011001010100001100000011",
    957 => "00111011001010010011101101111001",
    958 => "00111111100111001001111000110000",
    959 => "01011111010111001100110001111011",
    960 => "01010101101011001100100010100100",
    961 => "01010110100100101000111101011100",
    962 => "01001111000110110000110111100111",
    963 => "01011111001101001011110110001100",
    964 => "01011100011011110100010010100001",
    965 => "01010111101001001010110111100001",
    966 => "01010111001001111010101111110010",
    967 => "01001111100111001010000001101001",
    968 => "01011101000010110010010001110110",
    969 => "01011110101101000100001100110001",
    970 => "01011111011011110111001010101111",
    971 => "01011101101101000000111100110000",
    972 => "00101111000111011100011011111011",
    973 => "01010001101100101011111011001111",
    974 => "01000111011111111101110110011110",
    975 => "01001110011111111111010110101110",
    976 => "01001111101100110001101111100110",
    977 => "01000011101001110111011011001111",
    978 => "01001110100101111010010011001100",
    979 => "00110111101101000001011111001010",
    980 => "00101101001000111011100000111000",
    981 => "00111110101011101010011001010110",
    982 => "01011111000101010000110111101011",
    983 => "01000001101001011100001000011100",
    984 => "01001101101100000101110101110101",
    985 => "01010001101101001010110010110111",
    986 => "00111110111101000011000110111001",
    987 => "01000011010111001001010101011110",
    988 => "01001110111111111111010000100011",
    989 => "00111111101100110100111100110110",
    990 => "01011011101101000001111110111011",
    991 => "01010011101001110010010000111000",
    992 => "00110101010001010001110110010001",
    993 => "01011111011111101011010111111001",
    994 => "01010111001100011001001101001000",
    995 => "01010000100101011101110101000011",
    996 => "01011011101100011011001011010111",
    997 => "01001011101101001011000101010011",
    998 => "00110010100100101001110110100100",
    999 => "01010110111011110110101010010000");

  component fsqrt is
    port (A : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          Q : out std_logic_vector (31 downto 0));
  end component fsqrt;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (3 downto 0) of std_logic_vector (31 downto 0);
  signal cc : std_logic_vector (31 downto 0) := (others => '0');  
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0'); 
  signal Q_buff : std_logic_vector (7 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
  signal i_isRunning : std_logic := 'U';
  signal i_result : std_logic := '1';
begin  -- architecture fsqrt_tb

  i_fsqrt : fsqrt port map (s_a,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk,Q_buff) is
    variable ss : character;
    variable count : integer := 1;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      s_a <= a_lut (addr);
      cc <= ans_lut (addr);
      ccc <= cc ;

      if i_isRunning = '1' then  -- rising clock edge
        if ccc = c and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 1 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;

  end process ram_loop;

end architecture;
