library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity fabs_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity fabs_tb;

architecture testbench of fabs_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "10011111110110111101011010100110",
    1 => "01111101111100110101111100010101",
    2 => "11011111111111110111101010011100",
    3 => "10011111111101101111111111111000",
    4 => "11011111111111101011110101010011",
    5 => "11111101111111111000001101100010",
    6 => "01111111001111110000010010111000",
    7 => "10011111011111111001011100101100",
    8 => "01011101110000100011010111100111",
    9 => "00111011100101101010001000100000",
    10 => "11101111100111111000100010100010",
    11 => "11010001001111110100001110100000",
    12 => "11111001010111111001010111001001",
    13 => "01111100111011111111001101110101",
    14 => "01111010111111110011011110110001",
    15 => "11111110010111111110001001010010",
    16 => "11110111010110111110011111101110",
    17 => "11110101011001110100111111100010",
    18 => "11001011100111111000001000110101",
    19 => "01011111110111111111111000010001",
    20 => "00011110110011011001110110010101",
    21 => "01111110111011011000010011000010",
    22 => "01101111101111110101001001000011",
    23 => "11011011111111011110001110111111",
    24 => "01110111011111111111101111001111",
    25 => "11110110010111010101110000000101",
    26 => "11110111111011111101011011001010",
    27 => "11011110011111110101101010110000",
    28 => "11111110011011110101111000111101",
    29 => "01111101100111110001110011001010",
    30 => "00101110101110010100010010101111",
    31 => "11110111100100110010001011011010",
    32 => "10111111011011111010100111111010",
    33 => "11111101101111101010101010100110",
    34 => "00111111011110001010101011010101",
    35 => "01111101111011000011001001111101",
    36 => "10001111110101011110101000010001",
    37 => "01011100111110110101111110100110",
    38 => "10111111101011111111010100110000",
    39 => "11111011111111110001111101001100",
    40 => "00011011111111111001011000111010",
    41 => "11110111010001010000110001011110",
    42 => "01110011011111100100110001000101",
    43 => "01101111011000001011011110111101",
    44 => "01110011101111111110010110011111",
    45 => "01010111110011100001010000101111",
    46 => "11111110111111110000100111000011",
    47 => "10111101111111010100001110000010",
    48 => "11111001010111001110100110000100",
    49 => "01101110101011011111101011000000",
    50 => "01111011011101111010011000100001",
    51 => "11111111011111111010011110011010",
    52 => "11110110111001110001011000010001",
    53 => "11000011101110110110011101001100",
    54 => "11111101100001110100000011100011",
    55 => "01001111010011111100111101000000",
    56 => "01101110011010111001111001001111",
    57 => "11001011111011111000101010100101",
    58 => "10111110110111111100101000000000",
    59 => "11010011111101111100100110110101",
    60 => "01011111101111010101110110101011",
    61 => "01111011111110011000100001011100",
    62 => "01111101111000101000001100110111",
    63 => "01111101111111110010010000111001",
    64 => "11001011011111111011110010001000",
    65 => "01100101001110111101100001011101",
    66 => "11111110111111100110010110101100",
    67 => "11011110111111000010101100001001",
    68 => "01111011111111111011000111111000",
    69 => "10010101001110001100101001111110",
    70 => "01111111001111111011100100101110",
    71 => "01111111011011111110001101010000",
    72 => "10111111011111101101101101101100",
    73 => "10110101001001101100011000111000",
    74 => "01110111111001111000000100010100",
    75 => "01011011011100111011001001011010",
    76 => "00110101111111110110111111001101",
    77 => "11111110000101110111101101010000",
    78 => "00110111110111111011001110001001",
    79 => "11101011111011110101111001100001",
    80 => "11101110100111011001101111111100",
    81 => "11001111111111110111101001010101",
    82 => "00101101010011011001000100000101",
    83 => "01011011100011110011001011110010",
    84 => "11111101111000101010110110000110",
    85 => "01111010110011011101011010001011",
    86 => "10111111111111010100001110011101",
    87 => "00111111010011100111000110100111",
    88 => "11101110010001101100010000101100",
    89 => "01111110111101110101101111000011",
    90 => "11011011110111101111000110110000",
    91 => "01101111010100011010110000010111",
    92 => "01011111111011010101111110010111",
    93 => "11111101111110011010010011011010",
    94 => "01011100110101111110101110000111",
    95 => "01110101110111001000001000000101",
    96 => "00111011110111110000011111011011",
    97 => "00111110110011111001001000101001",
    98 => "01010101001110110010011011101101",
    99 => "01101111101010111000100111110011",
    100 => "01101110111001011000100110010101",
    101 => "01101111111101110011001101111011",
    102 => "11101111011111110100111001100001",
    103 => "01011110111101111100010001000111",
    104 => "01111110010111110101101011001111",
    105 => "11111010011111101010110100010011",
    106 => "01010011111011011100111111111111",
    107 => "11111011111001110111100001011110",
    108 => "11111110011101111001001011000011",
    109 => "10011110101111110010000101100010",
    110 => "01111011111110101101010101101100",
    111 => "11111100110110011111001100111011",
    112 => "01111101101111101100000100010010",
    113 => "11111011000011110110011011100100",
    114 => "11110011011110010111100011001001",
    115 => "11111110110101010010011000101000",
    116 => "01111110100110010011111000111010",
    117 => "00010110100010110011101110000011",
    118 => "10110110010100101011010010011011",
    119 => "01100111101111100111001011100000",
    120 => "01010010110111110101000010111000",
    121 => "11011001001111111011001110011011",
    122 => "01100111011111111111111001100101",
    123 => "00111111111101111100001101111001",
    124 => "11110010111011111110000011111101",
    125 => "11111110011011011101001101010010",
    126 => "11110110100111110100110011100000",
    127 => "00011111111100101011001011000010",
    128 => "01011011111101110100001110111100",
    129 => "10111100101111111100110111111001",
    130 => "11111110011110010000101000100000",
    131 => "01111011011110110110100011001010",
    132 => "10111101110011110110100010101011",
    133 => "00011111011011100100101011011100",
    134 => "11101111010111110111111011110101",
    135 => "00111111111101010000000010011011",
    136 => "01011111111111100111100011101111",
    137 => "01011011111011100001111011000111",
    138 => "11111011111111111110100011001100",
    139 => "00111111111011010001000001010101",
    140 => "11100111110111111011100010100111",
    141 => "11111100111001110100001110011110",
    142 => "00010001111110101101110010111110",
    143 => "11100110110111111011100011101001",
    144 => "00110101101111110000010110111001",
    145 => "01111110111111110010111100111010",
    146 => "01111110010111101100011000000000",
    147 => "01110110101111111000101110101011",
    148 => "01011110111011000011011111010011",
    149 => "01111110011111111000101111110110",
    150 => "11101110111110110011110100110000",
    151 => "11110111011111110011011101101111",
    152 => "01011111001111111111100001001001",
    153 => "11100011100111010001000000001011",
    154 => "01110111011111110100100001010000",
    155 => "00111011111111000001011011000001",
    156 => "01011110111111111110001101111000",
    157 => "11010010001101101111110101011011",
    158 => "01111011101100111010011100010101",
    159 => "11011111010111111101011111110111",
    160 => "10011101111101111110000000010101",
    161 => "01101011110010000101000001100110",
    162 => "10001010011110011001111010010110",
    163 => "01101011101111110111011001100000",
    164 => "11110011100101011100000010100111",
    165 => "11111011011111100000101011101111",
    166 => "01011011111111000110100110110000",
    167 => "01111011111111000100111001001101",
    168 => "11111111010111111001101000011100",
    169 => "01111101101101111001011110010101",
    170 => "10011100111100110101010101101110",
    171 => "11101001111111110011110111001011",
    172 => "11111110111010110100101100110101",
    173 => "00110111111111110011001100010110",
    174 => "00001011100101111100000100100100",
    175 => "01011111101111110111111011101100",
    176 => "11110111111111011001001111001111",
    177 => "01111101111101101000101001000111",
    178 => "11110101101101111010100011011110",
    179 => "10111011110111101001100001101111",
    180 => "01111110101111011000110001001010",
    181 => "00101111111001110011000101110111",
    182 => "11111101011111011010001111111011",
    183 => "11110001110101110101110111111110",
    184 => "10101011011101111000111010011111",
    185 => "11100001101111011100011010100111",
    186 => "11111011110101111100110001100000",
    187 => "10011111100001011101010011100001",
    188 => "01011011110111111000110101101101",
    189 => "00110011001111101110110101000000",
    190 => "11110111111110010111010110110010",
    191 => "11000011101111110000110010111110",
    192 => "11100111011011110000010010000111",
    193 => "10011000110111110101110100011001",
    194 => "10001110101100010010000111101011",
    195 => "11111101111101111011011100111001",
    196 => "01111011111111010101011110011110",
    197 => "10111101111111010110011011110000",
    198 => "11111101100111110011110011111011",
    199 => "00001011111111110101111011001111",
    200 => "00111011101110001011011101000100",
    201 => "11101101111011111000010101111001",
    202 => "00011010111111101011100010110101",
    203 => "10111111111101111101111111110100",
    204 => "01111011101011110011010000100010",
    205 => "10101101111111110001110101111100",
    206 => "01101010011111110001101100001000",
    207 => "11101011011011111100111101101001",
    208 => "11110001011101111011000001100001",
    209 => "01101111110111100101011110111110",
    210 => "10111111010111101000101100001010",
    211 => "11110001111110101100001011001111",
    212 => "11010111111010011110011110001001",
    213 => "10011111111011110000001101101100",
    214 => "11011110111101011110111011111000",
    215 => "01111010111010111001101111001011",
    216 => "11001111111111110100110110100010",
    217 => "01111111001111110011001111110111",
    218 => "01101110111111110111100111000001",
    219 => "11100111111101111001010101011001",
    220 => "01111110110011100110111010001110",
    221 => "00111111111111001010111100000011",
    222 => "01110110110010110101011000010110",
    223 => "11100111111011111000011010001010",
    224 => "01101101111111111011011000011110",
    225 => "00011111100111111101001100011011",
    226 => "10111010111011010100100100100011",
    227 => "01011110111111111101111011011110",
    228 => "11001101111111100101100101110011",
    229 => "10110111011101111101010101110100",
    230 => "01110011111111110111010110000011",
    231 => "11011111101111111000111101001111",
    232 => "11100111010101110100000100101100",
    233 => "11111110111111110010111001000100",
    234 => "11001111111111110001001001000101",
    235 => "10110000110101111010000011000011",
    236 => "01001111110111100010100001100000",
    237 => "01111111011101101001111111000011",
    238 => "01101111111011100101011010001000",
    239 => "00101111101111110101111110010111",
    240 => "01111010101100110110111110100111",
    241 => "11111011110010110010011110111100",
    242 => "01011111101110111110110101011000",
    243 => "01110110110110110000010101011010",
    244 => "11011010110111111101010001110001",
    245 => "01001011111101011100101100110010",
    246 => "01011010110111110100110000001110",
    247 => "11011101001111110000110100011010",
    248 => "00111011110111100001110111000111",
    249 => "00110001110111100100100000101001",
    250 => "11111000111111011111111011111100",
    251 => "01110111110111001011000011011111",
    252 => "01011010111000110011100010110011",
    253 => "10111111011110111010010111010010",
    254 => "01010101111011110111011011110001",
    255 => "11110111101110111001101111100001",
    256 => "11100111100111110011100000011101",
    257 => "00101101011101111001111101100011",
    258 => "10100110101111101100101000111000",
    259 => "10111110111110100110110001000000",
    260 => "01110111111101100111111110001101",
    261 => "11101011101110111110100010011111",
    262 => "11111101111110011001000111110011",
    263 => "10111111111111100101100011010110",
    264 => "00110010011101101101111111000110",
    265 => "11111101101101111000100111101100",
    266 => "11110110100111110101011101110000",
    267 => "11111111010101101110000101001000",
    268 => "01011000001111110101000111011010",
    269 => "11111101101111110000001010101100",
    270 => "11111111001101011011000101011000",
    271 => "01111011111110010110000000111110",
    272 => "11011110111111111000001011110011",
    273 => "01010010100100110001101000111011",
    274 => "01100011110110100000001111110000",
    275 => "11110111111100111100111000011100",
    276 => "00100110111111111111100010010011",
    277 => "01111111011100111100011111110010",
    278 => "01110111110111100101100110111111",
    279 => "11110001101011111011011000001001",
    280 => "11010111111100010001010001111101",
    281 => "01111111010111111010111001110010",
    282 => "11110001101111101110111110001011",
    283 => "00111110010111010101010000010010",
    284 => "00110101011010101110101111101000",
    285 => "01001101111111100000110010010010",
    286 => "11001111101011101000000011111011",
    287 => "11111011111101100001100010100101",
    288 => "00111100101101111001001000000110",
    289 => "01101010111110101001111000010000",
    290 => "10010110101011001011001001111001",
    291 => "11111011001111111000011100010101",
    292 => "01001111010101111100000001001111",
    293 => "01011110011111110001110101111010",
    294 => "11110111111001111010000011100101",
    295 => "10110101111101111100101100111110",
    296 => "01111010011111110001101110111001",
    297 => "01101111111010110010101011001111",
    298 => "01010111111101111000100010111100",
    299 => "10010111111011110111010100110101",
    300 => "11111110101110110110001011011101",
    301 => "11110111110110111001000101100111",
    302 => "01001111101111010001011011111110",
    303 => "10110110011110110100001010100111",
    304 => "01101111001001011110110100011010",
    305 => "11001111111111111010000001111010",
    306 => "01101011101111010011001110100100",
    307 => "01011111100110101110010101101001",
    308 => "01011001101111101111100011011000",
    309 => "10100011101101011100111011100101",
    310 => "01000110110111100010011011101111",
    311 => "10101111111111010001011011100100",
    312 => "00111011101111110011101001001011",
    313 => "11001111111100110000010101001111",
    314 => "11011111011011111111001010010100",
    315 => "00101001110100111111101100101011",
    316 => "11101111111011111110011111111000",
    317 => "00101111101100011010011110100101",
    318 => "11110111101111110100011110110010",
    319 => "11101100011011111000101011000001",
    320 => "11111110011001100010001010111110",
    321 => "01101110110111110101001111100110",
    322 => "00111001011011110101110011011111",
    323 => "01011101101101111100010100111001",
    324 => "11010100010111110100100110001000",
    325 => "01110010111101111101011101001100",
    326 => "01111110100111011111101001000100",
    327 => "01111100011111101101111000110111",
    328 => "11011101011010101001110011111011",
    329 => "10100111111101000010011000010000",
    330 => "11101101111101111001101010101001",
    331 => "11101011111111111010111110010100",
    332 => "01111010111111010110001001110101",
    333 => "10111101101101001100101010001001",
    334 => "01111110111011111111100010111011",
    335 => "01110111101111101110101101010011",
    336 => "10111000101111010101011110111110",
    337 => "11101001110011111010101101010010",
    338 => "10001111111111110100010010101011",
    339 => "01111100111111110001000110111110",
    340 => "00011100010010110111000011001111",
    341 => "10011110111111110010111101101001",
    342 => "01011111111010000000101110010110",
    343 => "11111100110110111011011100110110",
    344 => "11011111011011111110011100000011",
    345 => "11000111101011000010110110000110",
    346 => "11111101000111111010101011111101",
    347 => "01001101011110110110010000001000",
    348 => "00101111111100110001011101101111",
    349 => "00011011101011111001001010100110",
    350 => "01111101111111110100110100000000",
    351 => "10101101111111110110010111000101",
    352 => "00011111101101110010111010000111",
    353 => "01111011111100110100011000000101",
    354 => "01011111111101111001001110110110",
    355 => "00110100111011011001000000010111",
    356 => "10111111100001010110001111000110",
    357 => "01101111010111011001111100111101",
    358 => "01110111011111001100110100100000",
    359 => "10110110001000110001011111101110",
    360 => "01000111011111010011001110111011",
    361 => "10111101111111000010001010001110",
    362 => "00111011111111101110110000101010",
    363 => "00110111011010100100101000101001",
    364 => "11101111111011101111110011001011",
    365 => "00111111010100101011101000101001",
    366 => "00101110111011111100000100000110",
    367 => "00111110101111110101011111110010",
    368 => "10111111101110010101100101000001",
    369 => "11111010011111101110111000011011",
    370 => "10111111101111010010101100010101",
    371 => "01001011111110110100111011110010",
    372 => "10010110101011110110111101011111",
    373 => "11101101101011111000100001111000",
    374 => "10111111001101100110000101100101",
    375 => "01000111011110101110010100000100",
    376 => "01101111111011011100110001100001",
    377 => "11001001001111100001110011011100",
    378 => "11110111111101101101111100011100",
    379 => "11111101011011101111010001111110",
    380 => "10010011010100101101011100110101",
    381 => "01111111001111111111010011011110",
    382 => "01001110011111111100000110011110",
    383 => "10101111101110111110101011100000",
    384 => "00110111111111010100011010011101",
    385 => "10011111101100000110101011110101",
    386 => "11111010010101010101100011111000",
    387 => "11110111011101100001100000111101",
    388 => "01111101101110110111111110000100",
    389 => "10111110111011001000110001110111",
    390 => "01111001111111111100011100110011",
    391 => "10111111101101011100010111111110",
    392 => "11111010110110111010000010101001",
    393 => "01011101101111101011100111100001",
    394 => "10010111111101110001111111100111",
    395 => "00110111110101011110010001000000",
    396 => "10110111111111101100000000111101",
    397 => "10101011111111010110001011100100",
    398 => "11000110100011011100000100010010",
    399 => "00011111101010110011111100010001",
    400 => "01010111111011111001101011100010",
    401 => "01111010011111111111101101111011",
    402 => "10111111111111111101000011110010",
    403 => "10011101111111111101100011110011",
    404 => "10011110111111111111100101101110",
    405 => "10011011100111110010101110111001",
    406 => "10001011011111011000000111001101",
    407 => "01111011111011100001100111011100",
    408 => "01111011110110111101100110110111",
    409 => "11111101111111111100110011000100",
    410 => "11101101000101110100111010001000",
    411 => "10111011011111010110001111010110",
    412 => "11111001111111100011100000011111",
    413 => "11111011011111110101101011101101",
    414 => "00011110110111110001001100111100",
    415 => "00101110111111111111000101001110",
    416 => "11101110110010010010111101000101",
    417 => "00001111101111011001011010101010",
    418 => "10010101100110110101101001100101",
    419 => "10000110101111101010011100101010",
    420 => "00111010111111110010101000101111",
    421 => "01101101111011110000111010010111",
    422 => "11111010010011100110010010100101",
    423 => "01110001111011010111110111001110",
    424 => "11101111111111101010011001000101",
    425 => "01011111101110111011111001101011",
    426 => "01000010111110100111001010101111",
    427 => "01110111111111010101001001100011",
    428 => "11110101101110010001000110110000",
    429 => "10111111110110100010011000111101",
    430 => "11111100101101111000100111100000",
    431 => "00111101100011110011100001110011",
    432 => "01111110111111110000011011000000",
    433 => "00010101110111110101101000000010",
    434 => "00111101111111101111110110100101",
    435 => "11100011111111101111000000010001",
    436 => "11101110111111011111000011010011",
    437 => "01110111100011111010010100000110",
    438 => "10010100111111100100011101000101",
    439 => "11111101111101111010111100010100",
    440 => "01100101011111111001011110111010",
    441 => "10111001111010110001110111110001",
    442 => "01101111011111111000001100011111",
    443 => "01011111000011110101000111000100",
    444 => "11001110101101111100010011010000",
    445 => "11101011111100010011111000001011",
    446 => "11011100111111011110110011011010",
    447 => "10111111101111101110000011100111",
    448 => "11011110101111100101011010110101",
    449 => "01100110111011111011100000000100",
    450 => "10101100111111111000001001110111",
    451 => "01111101111111111111010101000011",
    452 => "11011111110010110001011101101101",
    453 => "01011111101110111010001000001100",
    454 => "01110001011101010010111100001100",
    455 => "11111110111101100001100010100111",
    456 => "00110110100111000101001010011000",
    457 => "11100011111101000111101011000111",
    458 => "00111010111100110100110000101100",
    459 => "01111101101011110000101100101000",
    460 => "11111110101111111011100011010000",
    461 => "00001111100001101100110010001110",
    462 => "11100101100110111100101010011100",
    463 => "01111101001100110101011001001101",
    464 => "01101111111110000010110101101010",
    465 => "01111101110101110111110110010000",
    466 => "01110100111111101010001110001001",
    467 => "11111101001111110111000010111101",
    468 => "11000111110101111101101110101100",
    469 => "01101011111111111111001011001001",
    470 => "01101101101101111001100100001110",
    471 => "01111011111111100000110111010001",
    472 => "01111011111111111010110100100111",
    473 => "11111101011011111001110010001001",
    474 => "01110101010111011001001100000011",
    475 => "01101110111110110110010011011111",
    476 => "11111011011011101110010000100011",
    477 => "00011011111111111011110000001110",
    478 => "00111111111111100000011010111101",
    479 => "11111100111101110101011001100100",
    480 => "11111001111111100101100100111010",
    481 => "11111101111110110000000101111110",
    482 => "11111101111110111011011000011110",
    483 => "11111110111001111000110101001110",
    484 => "00110110111111000010100100000111",
    485 => "11100111101111111010001000100010",
    486 => "01111110111011111001000011010101",
    487 => "00111111111111000111101111101110",
    488 => "01111101110111111001010000000100",
    489 => "11111011111101101000001101101001",
    490 => "01101111101111011000111101001000",
    491 => "01101011111101101011010000010000",
    492 => "11111110110111010111100100011010",
    493 => "11111111011111111000010011110100",
    494 => "11011111011111111010011101100101",
    495 => "10101110111110111100100101101100",
    496 => "01110101011111111000011000001101",
    497 => "10111111101111010010100001110010",
    498 => "11111101111111111110010111101100",
    499 => "01111110110000010000001010001001",
    500 => "11110111111110101001101010011001",
    501 => "01111110011111111100100110000110",
    502 => "01111101110111111000010110001111",
    503 => "11111110101110010111100101100100",
    504 => "11111110110110110011100001100100",
    505 => "10010111101101001101110010000111",
    506 => "10101101111011111000100010101100",
    507 => "10100111111110110111111001111011",
    508 => "10110101100001100001001111100111",
    509 => "01110001101111110001101001111100",
    510 => "10111101111101111111111101111100",
    511 => "11011110011100010010000100101000",
    512 => "11101111101011101101001100011000",
    513 => "01011101111001111100110001001110",
    514 => "01100111111111110110100001000101",
    515 => "11110100101010100101011101010000",
    516 => "01111101011110010100010000001011",
    517 => "01110011111110101000000001110011",
    518 => "01001001101001011011110100001100",
    519 => "11010110101010111010010101000001",
    520 => "01011111111111000001011111011010",
    521 => "11011101111111010001001110111100",
    522 => "11011110001111000111010101011001",
    523 => "10011011010011100111100101100011",
    524 => "11010111111001010001001100111100",
    525 => "01011111101111101101100111000110",
    526 => "11111110111111110100100011110110",
    527 => "01111100110111111011000011111001",
    528 => "01101101111011110111010010110110",
    529 => "11111101100001101100001011111010",
    530 => "00010111011001111110111010001100",
    531 => "01101111111111111111000101111110",
    532 => "10101110110011100010011110011000",
    533 => "11101110111110110111100000011111",
    534 => "11001111111111011000001010110101",
    535 => "10011110111100110010110000111101",
    536 => "10111001101101100110010110100010",
    537 => "11111111001001110010100010101010",
    538 => "00111011111011100010101011010111",
    539 => "00000101100111010111001011100101",
    540 => "10111011110111110100111010011111",
    541 => "11101111111011111101011111101010",
    542 => "01111100111001100111110011100000",
    543 => "01110011110101010001100010100110",
    544 => "01101110011111010100011011100000",
    545 => "01101111011111101001000010010101",
    546 => "01001000101111101011100010101111",
    547 => "00111011111001110011101101010001",
    548 => "01100111101111111001100010101110",
    549 => "11111110010100001101000111010111",
    550 => "11111010101011010000100100100101",
    551 => "01111011111111001101110101010101",
    552 => "01110011011110110011011001100111",
    553 => "10000101011001100011100010011001",
    554 => "01111100101111010000110000010110",
    555 => "11111110111110101000010010011111",
    556 => "01110111111111110001110101001100",
    557 => "01111110011101010011000010100000",
    558 => "01011001010011110100000101011010",
    559 => "11101000101110110111000111101011",
    560 => "00011011110101000101001101101100",
    561 => "00101100000111111111011010110011",
    562 => "00111011000111110000101100110100",
    563 => "01011111110111111001100110010100",
    564 => "10111110111111111010001000110010",
    565 => "01111110010001101101011010110110",
    566 => "01111111011011111100111111000011",
    567 => "01011011111101010100011101110100",
    568 => "01111101111011001011111111011010",
    569 => "11110010111110100101010101100101",
    570 => "11111110111111111011010100010101",
    571 => "01101111001111100011100111000001",
    572 => "11111101011011110001111011111010",
    573 => "00111111111011100010100110000000",
    574 => "01110100101101011001100101001001",
    575 => "11101100111110110100011110110011",
    576 => "11110111010111111101100010010111",
    577 => "01111010111111101111101000100001",
    578 => "01101111111111011000010000000000",
    579 => "01111010111111111111101001010010",
    580 => "11111111001111010101100000111001",
    581 => "01110111110110010111101101100101",
    582 => "11111000111010100001011000111010",
    583 => "11111011010011110101011001000011",
    584 => "11010010000001000110011110001010",
    585 => "10100110110011011111001001010000",
    586 => "01011111110100110001110100110010",
    587 => "11111110111110111001110000110010",
    588 => "11111011111001010101000010000101",
    589 => "01111111010111011001011101000100",
    590 => "11011111011111111100010100101100",
    591 => "01001011111011111010001111100111",
    592 => "11011110101111011001111101011111",
    593 => "11110111110111101010001111100011",
    594 => "01101101111011010110100001001110",
    595 => "01001111101111000001111100011000",
    596 => "11111010111111111011111101100011",
    597 => "11110101111111110111010000000101",
    598 => "11011111010111110110101101001000",
    599 => "11110110110101101010000011101101",
    600 => "11111111001111010101101001001100",
    601 => "01110111011111100101100101010111",
    602 => "11111101110011011010111100001101",
    603 => "11011101101111111101100101101111",
    604 => "11110110000101111110011111001000",
    605 => "11111011101111000110101011010000",
    606 => "11011111000111111110110110011011",
    607 => "00001100101101111001100110010101",
    608 => "01011010111110011110000101011010",
    609 => "01110111111111111010011100110001",
    610 => "01010110111111110010111010010110",
    611 => "11011111101100110001111110100111",
    612 => "01111011111101001110010101001100",
    613 => "00111110101011110110001011000000",
    614 => "00010011110011101111000101110010",
    615 => "00111111011011010011010000101101",
    616 => "00111101111111010001000101100001",
    617 => "00111111111111011110010010101010",
    618 => "00111011111011111010110000110111",
    619 => "10110101100011110000011010101000",
    620 => "00011110111011110001111110101100",
    621 => "11111001011001010100010010010110",
    622 => "01110111111110010010101110011110",
    623 => "11011010110110010001001000111010",
    624 => "01001100110110110111101101010000",
    625 => "11011111111111111110010101001010",
    626 => "11001110110111100001000001010100",
    627 => "01110111101101110001010011101011",
    628 => "01001111110111100000100100111010",
    629 => "01111101111101111000010011100011",
    630 => "10010110110011010010010111001010",
    631 => "00001111011101100100101100000011",
    632 => "11110111101111101101000001010101",
    633 => "11110111111111110100010111000001",
    634 => "11111010111011110100100001110101",
    635 => "10011101010011111001010111111100",
    636 => "11100001110111110110010000101000",
    637 => "01110111111111111011001011111011",
    638 => "01101110110111111001010001101011",
    639 => "01111011101111111011011100110011",
    640 => "11100111110011011100100101000011",
    641 => "11111110111011110100010001001011",
    642 => "01101111110101010011101010011101",
    643 => "01001010111111101000101011101100",
    644 => "11010111111011110101010111000100",
    645 => "00111110001110010001010011001010",
    646 => "01011010101111101100110100101010",
    647 => "01111111011001011111110100010110",
    648 => "01001111110010111101000110011101",
    649 => "01101111100111100000001101001011",
    650 => "01100111011101111101001010010110",
    651 => "11111101101111010010100100110101",
    652 => "11111101101001111101110111010101",
    653 => "10011101001111111011001111011101",
    654 => "01111101101000100011011101010101",
    655 => "11010111011011100101101101001110",
    656 => "01110110101100110101011010101110",
    657 => "11101100011110110100101000110001",
    658 => "01011110111111000010101000000010",
    659 => "11110111101111101101001010001011",
    660 => "10011111001001010100111110010000",
    661 => "01011011111111110001010100101100",
    662 => "11101111111001111111001010111111",
    663 => "00011011111111101011101001001110",
    664 => "10011010001111010110110101010011",
    665 => "01101001011111001101100110010100",
    666 => "01010001111011010010110100101101",
    667 => "10101001111111101001111001010000",
    668 => "11111011100111111000110010001010",
    669 => "01010101111101010010000011101100",
    670 => "10011111111010111010100111000010",
    671 => "11111110110111111110001010100111",
    672 => "11011100111111111100101011110000",
    673 => "01011011100011011100011000111000",
    674 => "11011011111111000010011101010101",
    675 => "01011010010101000110110101011100",
    676 => "01110111111110111100001100100110",
    677 => "01110100011111010011011000001001",
    678 => "01001111110111011011111111001111",
    679 => "11111110111111110101000110101010",
    680 => "10111111111100010111011010111010",
    681 => "10111111101001101110100110011001",
    682 => "00110111111100110000001011000001",
    683 => "10101111111011110000111101000000",
    684 => "00110011110111001010011010111111",
    685 => "11011101011011101000000001001000",
    686 => "01101011001110100010100111100011",
    687 => "11110000000110110010010110010110",
    688 => "01101100111111110110010110111001",
    689 => "11010111100101111100101101111111",
    690 => "10001110111011110110011011111111",
    691 => "10111101001011001111101011000001",
    692 => "10111011111110001011111100011110",
    693 => "00010100111111011010110010100110",
    694 => "11001111101011011010011110001100",
    695 => "01011111011101100000000011000011",
    696 => "11111111011111100111101000111110",
    697 => "01111110111111111011010111101100",
    698 => "11100101111011000000110101110000",
    699 => "10110101111011110010100110000010",
    700 => "10111101111110101111100001111000",
    701 => "00100110011111110011110110010101",
    702 => "01101111001111111111010100000011",
    703 => "01111110111111100001001001110110",
    704 => "11111101111111111011000000010110",
    705 => "00111111111101110010110111010010",
    706 => "00111111111100110110110010011010",
    707 => "01101011101111011011010000011110",
    708 => "01110011110101001110001100100011",
    709 => "10111011101011110011110010000001",
    710 => "00111111011011100010110111110001",
    711 => "10101101011011111010100011110101",
    712 => "01111110111010010010011110100000",
    713 => "01111101110100100010010100101110",
    714 => "01011110110001011110100100111111",
    715 => "00100111110101011111100001111011",
    716 => "11101101011111100011111011100000",
    717 => "00111110011111110100100000111011",
    718 => "01110110010111110010111101001011",
    719 => "10111011111101110101000100101101",
    720 => "01000101110010111001111010100001",
    721 => "11000011110011011100011110011110",
    722 => "00001111000111110110011000010000",
    723 => "10110110010100010000110001110100",
    724 => "11110111011011110100000101100011",
    725 => "01111001101111110011110000110001",
    726 => "01111111010111110001010001001011",
    727 => "00111101111111001001111000010100",
    728 => "10101111010111111011000000010000",
    729 => "10111000101111110101010011011110",
    730 => "10110111111111111010111000101000",
    731 => "01111101001011011001011000001010",
    732 => "11011111011111011110010100010101",
    733 => "00011100011001000111001001000000",
    734 => "11011111011011110101010001010011",
    735 => "01110111111111101100100010111000",
    736 => "00111110111011110111010010111000",
    737 => "11110011101011010111110000000011",
    738 => "10111111011101111100001011001010",
    739 => "11111110111111110011011010010110",
    740 => "01011110111001110010011001101001",
    741 => "11101101111111110110000001011010",
    742 => "01010100011010111000001100111001",
    743 => "11011000000101110100101111010001",
    744 => "11111101111110111011100011110111",
    745 => "01011111111110110110101111010110",
    746 => "01011011111110110011001000100010",
    747 => "11100110111110100010110101000111",
    748 => "11101111110111100110010101001011",
    749 => "01010101111100010110011111001111",
    750 => "11101101010111111000110101110101",
    751 => "00011101011111100101111101010000",
    752 => "00110110010110100110101001110011",
    753 => "10101011001011111100011011011110",
    754 => "11101101011011000010000100010101",
    755 => "11101101111100001110101111101010",
    756 => "11111101111111101001000111011011",
    757 => "01101110111100110100011100111011",
    758 => "10110011011111011111011110010000",
    759 => "01101011101110111001100111010011",
    760 => "11010111001111100000001111111100",
    761 => "11111111011011100111111011011001",
    762 => "01101101010111100110011001101100",
    763 => "11011111111111011010011010001001",
    764 => "01010000111111010001010111000111",
    765 => "00101000111111011011001000000101",
    766 => "10111111111011111100100111101101",
    767 => "01011100111110010000110100010010",
    768 => "01111101111011110111100101001001",
    769 => "01111101111110110110011100001010",
    770 => "01111011111111110000011101011110",
    771 => "01101011011110111001101010001100",
    772 => "01101101111001111100011111111000",
    773 => "00010111111011100111010010100010",
    774 => "11110111011110111001111010000101",
    775 => "01000110111110111100110111101111",
    776 => "01111111011110001111111111001001",
    777 => "01110111101101111100101010101111",
    778 => "10111010111111111000010101110100",
    779 => "00110111011110011111001000110110",
    780 => "01110111110110011101010101101000",
    781 => "11111011111111110011011111010110",
    782 => "10110011111010110110001000001000",
    783 => "11001111111111110011011011001000",
    784 => "00111110011011100010000111111001",
    785 => "10111101111011111100100111110000",
    786 => "10011101111010010100100110000001",
    787 => "11010011111111101010001010010100",
    788 => "01110000100110111011000110011110",
    789 => "10111011111111111110010011111011",
    790 => "01111111011111111100011011111000",
    791 => "11111101111011100100010111010011",
    792 => "01010011010011111010000111101000",
    793 => "11101101001010110100011100010111",
    794 => "10111011001111010101100111001011",
    795 => "10111110110110110101111001001000",
    796 => "11000010111101010111001000110010",
    797 => "00111101101111111100111010111001",
    798 => "01011011111110110011110011000111",
    799 => "01111101111111111100111000001010",
    800 => "01111000110111111101011001011101",
    801 => "11101110101111111110000100100010",
    802 => "11110111110111110011100101100011",
    803 => "00101101011111111000000110000100",
    804 => "11010111111110000011000010001101",
    805 => "11011011111101101011100110001001",
    806 => "01111110110111111100100010011111",
    807 => "00101111111101110100100111000110",
    808 => "10101011100111011101110000000010",
    809 => "00111111010011111011100011010110",
    810 => "00111011111111010011010000100100",
    811 => "00000011110111111011101010001100",
    812 => "11111111010111110110011100101011",
    813 => "00111101111101100001101100011000",
    814 => "11111011011111100101100101000000",
    815 => "10001110111101110111100101110001",
    816 => "10110010110111000110110100010001",
    817 => "01111101101110111011001100101111",
    818 => "01101100101110111011010111101110",
    819 => "01111110110011110101000000011001",
    820 => "01111111011111110011110101110001",
    821 => "01111001100101111011000111100000",
    822 => "01111100011011110111001000100011",
    823 => "11011001011011110111010001110011",
    824 => "11111101111111110000111010000100",
    825 => "10111100011111111000000100000010",
    826 => "11111110011111110011101111011001",
    827 => "11101101111111110011101101010001",
    828 => "11011101011001101010110101001000",
    829 => "01111100011101111001011110000001",
    830 => "01011101011011110000011000001001",
    831 => "01010110011000101100110100110000",
    832 => "01101110111000111100101111111100",
    833 => "01011111011111111111000000000010",
    834 => "01111101111111111110000001011000",
    835 => "11011011111110001010000101011001",
    836 => "01110011011111101001111100001000",
    837 => "01111011111111011111111010100100",
    838 => "01101010111111111110110011001011",
    839 => "11111011011011111010001100001000",
    840 => "01100101000110110001111101100011",
    841 => "01011011001111101010111110101001",
    842 => "11101110111111110001111001111101",
    843 => "11001111110001110000010000100111",
    844 => "01111011111110110010110000111101",
    845 => "10111101000110111100111110001100",
    846 => "01010010100110010000111101010011",
    847 => "10110011111011111110110100000001",
    848 => "10001101111110101101010011000001",
    849 => "11011011111111011100010000101001",
    850 => "10110101111101001001111110000110",
    851 => "01011111110111100011010111001001",
    852 => "01011101001011011010110001000011",
    853 => "01011011111111100110011010011000",
    854 => "10001101110111111011000001101000",
    855 => "10111111101111110100011011100110",
    856 => "11111011011101110101000011011011",
    857 => "01111101111111010101000000111000",
    858 => "01111011111100110011001110110001",
    859 => "01000011001111010111011010000101",
    860 => "11111001111111111110111001100011",
    861 => "01110010101011100011101111010111",
    862 => "11111011111111011100001101100100",
    863 => "11111011111111110010001110000000",
    864 => "11101111110000110001110111101011",
    865 => "11110100111101110100111001011001",
    866 => "01111010101101110000100110011001",
    867 => "01011110011101101011001101010001",
    868 => "00110011100111110010110011011101",
    869 => "01100011110111101101011110001100",
    870 => "01111110111101010011110011011010",
    871 => "00111011001111110110001111001100",
    872 => "00101110111110100010011011000110",
    873 => "01000111011000110010100011110100",
    874 => "11011111010101111101011001100101",
    875 => "00110110111111110011001000000010",
    876 => "11111101011001100100100111100011",
    877 => "01101101011011111110110110011010",
    878 => "00111110111111000011110100100110",
    879 => "01101000111101111001000000001001",
    880 => "11111101111011100011101110101101",
    881 => "11101111111111111101101101101101",
    882 => "00011000010010101111010000010110",
    883 => "11001111101100101111001010001001",
    884 => "01101111111100110110100011011001",
    885 => "11011111101101010001100110110011",
    886 => "01010010011110010101101010100000",
    887 => "10100011110111111111001100111101",
    888 => "11101111101001111000001001111101",
    889 => "10110100011111110101101011101011",
    890 => "10101100110111111101101111011111",
    891 => "11101101111111111010100111100101",
    892 => "10111111011111000001001000110001",
    893 => "01011111111110101101010100000000",
    894 => "01101101100010011101010101100100",
    895 => "01110001011111011011100000101110",
    896 => "11010111101110111111111010101100",
    897 => "11110110111110100000000000010000",
    898 => "11110011110111111001101111100110",
    899 => "00101110101111111011111001100101",
    900 => "11011010100111100010000111111100",
    901 => "11001101111010010001100010010010",
    902 => "10111111110011110000000000110001",
    903 => "01011011010111011000111001000011",
    904 => "01111110011011110100111110001110",
    905 => "11111111011100111111111111101011",
    906 => "01011111110111010011001110011101",
    907 => "01001111111111111001000111101011",
    908 => "01100111110111110110000101110101",
    909 => "01011101101110110110110110100110",
    910 => "01111110111100100111100001100000",
    911 => "01111110111100011010110100111111",
    912 => "01101001011101110101111100010101",
    913 => "01111111011110110110101100001010",
    914 => "10111111001001110100110111100100",
    915 => "00011111110011101111010110010010",
    916 => "00101111111111000000100110100100",
    917 => "01011111111101011110001111101001",
    918 => "01111010101011101010100100110011",
    919 => "01110100111111111101110001001111",
    920 => "00111111111011101111001000110100",
    921 => "11101100111111110111011011111011",
    922 => "11111111011101010001100010001001",
    923 => "10100111101110001110101101101110",
    924 => "01100111111011111111001000010011",
    925 => "10011111011100101111001010000010",
    926 => "01010011111101111101110001000000",
    927 => "01010111011110101110100001110111",
    928 => "01111111010110110110111100010001",
    929 => "01100111111011101101010001010001",
    930 => "11011101111111010101010110100011",
    931 => "00111001100011110111001011001000",
    932 => "01011111111111001110011111001011",
    933 => "01011110111111011010101110111001",
    934 => "10101011110010110001010010111101",
    935 => "00101110111110101011000110011011",
    936 => "00111000100111101001011111110101",
    937 => "11110101111111111000101100010001",
    938 => "01111110111001010000000100000110",
    939 => "11110111110110100011011010101110",
    940 => "01111110111111000111101011001000",
    941 => "11010111111010111011000100111111",
    942 => "00000111111010110100111001111110",
    943 => "11000011110111101011000000100000",
    944 => "11010111111010110100000001101111",
    945 => "11110110110000101110010010101001",
    946 => "10111110011111010111010000110001",
    947 => "00001100101101101111100011110010",
    948 => "11111100111010111011111011011011",
    949 => "11110111011100111111101010000011",
    950 => "11110111110101111011001011111011",
    951 => "01100101111011010001110010000100",
    952 => "11011111111111101000101101100001",
    953 => "11101111101110111100000001001100",
    954 => "01101011100011100111100001101110",
    955 => "10111001111111111001000011101011",
    956 => "01101110001111011010001101110010",
    957 => "11001110111110111010010100000110",
    958 => "00111101111111110110000000101101",
    959 => "01111111001111110001111001011111",
    960 => "11111101101110110010010101011101",
    961 => "11110011111010111101110100100011",
    962 => "11011111111011101001110100011100",
    963 => "01010111010111111101010101010101",
    964 => "00110111111110111001010101111111",
    965 => "01110111110110111000100100100101",
    966 => "01001111110111011100000100010101",
    967 => "01011100111111111100011101010111",
    968 => "00111111111001011101100111110000",
    969 => "01111011111111110010100000000010",
    970 => "11011111011111101111100010100011",
    971 => "11111101101110111101100100001001",
    972 => "01111001001101110101001110001111",
    973 => "01111101111011111011011011100001",
    974 => "11111110111111111001001001010110",
    975 => "01111111011111110100111100101001",
    976 => "11101110010011011011111001000001",
    977 => "11010111100101100100011100011111",
    978 => "11110101110111001000010101101111",
    979 => "01001111111101000010101101110011",
    980 => "11111100101010000010011110100111",
    981 => "11101110111111110001100011100000",
    982 => "01111111011101100010111011000100",
    983 => "01100111111001110101110110101100",
    984 => "00111111111101111111110001111010",
    985 => "01010000010111111100010100010001",
    986 => "01111011111110110110111111101100",
    987 => "01000010011000111100000111110111",
    988 => "00011001111010000101100000110010",
    989 => "01111111011110110111000110111011",
    990 => "10111111111111101111110101100101",
    991 => "00111101111001101010101000001001",
    992 => "00111111111110111010110001110011",
    993 => "11010111111111110000101110011110",
    994 => "01110111110101010011111000001100",
    995 => "01111110111111011100010001101110",
    996 => "11001101011111110010001001000100",
    997 => "10100111111010101111111001111000",
    998 => "11111011111110100111100001101111",
    999 => "01111101100110011101111000100000");

  constant ans_lut : lut := (
    0 => "00011111110110111101011010100110",
    1 => "01111101111100110101111100010101",
    2 => "01011111111111110111101010011100",
    3 => "00011111111101101111111111111000",
    4 => "01011111111111101011110101010011",
    5 => "01111101111111111000001101100010",
    6 => "01111111001111110000010010111000",
    7 => "00011111011111111001011100101100",
    8 => "01011101110000100011010111100111",
    9 => "00111011100101101010001000100000",
    10 => "01101111100111111000100010100010",
    11 => "01010001001111110100001110100000",
    12 => "01111001010111111001010111001001",
    13 => "01111100111011111111001101110101",
    14 => "01111010111111110011011110110001",
    15 => "01111110010111111110001001010010",
    16 => "01110111010110111110011111101110",
    17 => "01110101011001110100111111100010",
    18 => "01001011100111111000001000110101",
    19 => "01011111110111111111111000010001",
    20 => "00011110110011011001110110010101",
    21 => "01111110111011011000010011000010",
    22 => "01101111101111110101001001000011",
    23 => "01011011111111011110001110111111",
    24 => "01110111011111111111101111001111",
    25 => "01110110010111010101110000000101",
    26 => "01110111111011111101011011001010",
    27 => "01011110011111110101101010110000",
    28 => "01111110011011110101111000111101",
    29 => "01111101100111110001110011001010",
    30 => "00101110101110010100010010101111",
    31 => "01110111100100110010001011011010",
    32 => "00111111011011111010100111111010",
    33 => "01111101101111101010101010100110",
    34 => "00111111011110001010101011010101",
    35 => "01111101111011000011001001111101",
    36 => "00001111110101011110101000010001",
    37 => "01011100111110110101111110100110",
    38 => "00111111101011111111010100110000",
    39 => "01111011111111110001111101001100",
    40 => "00011011111111111001011000111010",
    41 => "01110111010001010000110001011110",
    42 => "01110011011111100100110001000101",
    43 => "01101111011000001011011110111101",
    44 => "01110011101111111110010110011111",
    45 => "01010111110011100001010000101111",
    46 => "01111110111111110000100111000011",
    47 => "00111101111111010100001110000010",
    48 => "01111001010111001110100110000100",
    49 => "01101110101011011111101011000000",
    50 => "01111011011101111010011000100001",
    51 => "01111111011111111010011110011010",
    52 => "01110110111001110001011000010001",
    53 => "01000011101110110110011101001100",
    54 => "01111101100001110100000011100011",
    55 => "01001111010011111100111101000000",
    56 => "01101110011010111001111001001111",
    57 => "01001011111011111000101010100101",
    58 => "00111110110111111100101000000000",
    59 => "01010011111101111100100110110101",
    60 => "01011111101111010101110110101011",
    61 => "01111011111110011000100001011100",
    62 => "01111101111000101000001100110111",
    63 => "01111101111111110010010000111001",
    64 => "01001011011111111011110010001000",
    65 => "01100101001110111101100001011101",
    66 => "01111110111111100110010110101100",
    67 => "01011110111111000010101100001001",
    68 => "01111011111111111011000111111000",
    69 => "00010101001110001100101001111110",
    70 => "01111111001111111011100100101110",
    71 => "01111111011011111110001101010000",
    72 => "00111111011111101101101101101100",
    73 => "00110101001001101100011000111000",
    74 => "01110111111001111000000100010100",
    75 => "01011011011100111011001001011010",
    76 => "00110101111111110110111111001101",
    77 => "01111110000101110111101101010000",
    78 => "00110111110111111011001110001001",
    79 => "01101011111011110101111001100001",
    80 => "01101110100111011001101111111100",
    81 => "01001111111111110111101001010101",
    82 => "00101101010011011001000100000101",
    83 => "01011011100011110011001011110010",
    84 => "01111101111000101010110110000110",
    85 => "01111010110011011101011010001011",
    86 => "00111111111111010100001110011101",
    87 => "00111111010011100111000110100111",
    88 => "01101110010001101100010000101100",
    89 => "01111110111101110101101111000011",
    90 => "01011011110111101111000110110000",
    91 => "01101111010100011010110000010111",
    92 => "01011111111011010101111110010111",
    93 => "01111101111110011010010011011010",
    94 => "01011100110101111110101110000111",
    95 => "01110101110111001000001000000101",
    96 => "00111011110111110000011111011011",
    97 => "00111110110011111001001000101001",
    98 => "01010101001110110010011011101101",
    99 => "01101111101010111000100111110011",
    100 => "01101110111001011000100110010101",
    101 => "01101111111101110011001101111011",
    102 => "01101111011111110100111001100001",
    103 => "01011110111101111100010001000111",
    104 => "01111110010111110101101011001111",
    105 => "01111010011111101010110100010011",
    106 => "01010011111011011100111111111111",
    107 => "01111011111001110111100001011110",
    108 => "01111110011101111001001011000011",
    109 => "00011110101111110010000101100010",
    110 => "01111011111110101101010101101100",
    111 => "01111100110110011111001100111011",
    112 => "01111101101111101100000100010010",
    113 => "01111011000011110110011011100100",
    114 => "01110011011110010111100011001001",
    115 => "01111110110101010010011000101000",
    116 => "01111110100110010011111000111010",
    117 => "00010110100010110011101110000011",
    118 => "00110110010100101011010010011011",
    119 => "01100111101111100111001011100000",
    120 => "01010010110111110101000010111000",
    121 => "01011001001111111011001110011011",
    122 => "01100111011111111111111001100101",
    123 => "00111111111101111100001101111001",
    124 => "01110010111011111110000011111101",
    125 => "01111110011011011101001101010010",
    126 => "01110110100111110100110011100000",
    127 => "00011111111100101011001011000010",
    128 => "01011011111101110100001110111100",
    129 => "00111100101111111100110111111001",
    130 => "01111110011110010000101000100000",
    131 => "01111011011110110110100011001010",
    132 => "00111101110011110110100010101011",
    133 => "00011111011011100100101011011100",
    134 => "01101111010111110111111011110101",
    135 => "00111111111101010000000010011011",
    136 => "01011111111111100111100011101111",
    137 => "01011011111011100001111011000111",
    138 => "01111011111111111110100011001100",
    139 => "00111111111011010001000001010101",
    140 => "01100111110111111011100010100111",
    141 => "01111100111001110100001110011110",
    142 => "00010001111110101101110010111110",
    143 => "01100110110111111011100011101001",
    144 => "00110101101111110000010110111001",
    145 => "01111110111111110010111100111010",
    146 => "01111110010111101100011000000000",
    147 => "01110110101111111000101110101011",
    148 => "01011110111011000011011111010011",
    149 => "01111110011111111000101111110110",
    150 => "01101110111110110011110100110000",
    151 => "01110111011111110011011101101111",
    152 => "01011111001111111111100001001001",
    153 => "01100011100111010001000000001011",
    154 => "01110111011111110100100001010000",
    155 => "00111011111111000001011011000001",
    156 => "01011110111111111110001101111000",
    157 => "01010010001101101111110101011011",
    158 => "01111011101100111010011100010101",
    159 => "01011111010111111101011111110111",
    160 => "00011101111101111110000000010101",
    161 => "01101011110010000101000001100110",
    162 => "00001010011110011001111010010110",
    163 => "01101011101111110111011001100000",
    164 => "01110011100101011100000010100111",
    165 => "01111011011111100000101011101111",
    166 => "01011011111111000110100110110000",
    167 => "01111011111111000100111001001101",
    168 => "01111111010111111001101000011100",
    169 => "01111101101101111001011110010101",
    170 => "00011100111100110101010101101110",
    171 => "01101001111111110011110111001011",
    172 => "01111110111010110100101100110101",
    173 => "00110111111111110011001100010110",
    174 => "00001011100101111100000100100100",
    175 => "01011111101111110111111011101100",
    176 => "01110111111111011001001111001111",
    177 => "01111101111101101000101001000111",
    178 => "01110101101101111010100011011110",
    179 => "00111011110111101001100001101111",
    180 => "01111110101111011000110001001010",
    181 => "00101111111001110011000101110111",
    182 => "01111101011111011010001111111011",
    183 => "01110001110101110101110111111110",
    184 => "00101011011101111000111010011111",
    185 => "01100001101111011100011010100111",
    186 => "01111011110101111100110001100000",
    187 => "00011111100001011101010011100001",
    188 => "01011011110111111000110101101101",
    189 => "00110011001111101110110101000000",
    190 => "01110111111110010111010110110010",
    191 => "01000011101111110000110010111110",
    192 => "01100111011011110000010010000111",
    193 => "00011000110111110101110100011001",
    194 => "00001110101100010010000111101011",
    195 => "01111101111101111011011100111001",
    196 => "01111011111111010101011110011110",
    197 => "00111101111111010110011011110000",
    198 => "01111101100111110011110011111011",
    199 => "00001011111111110101111011001111",
    200 => "00111011101110001011011101000100",
    201 => "01101101111011111000010101111001",
    202 => "00011010111111101011100010110101",
    203 => "00111111111101111101111111110100",
    204 => "01111011101011110011010000100010",
    205 => "00101101111111110001110101111100",
    206 => "01101010011111110001101100001000",
    207 => "01101011011011111100111101101001",
    208 => "01110001011101111011000001100001",
    209 => "01101111110111100101011110111110",
    210 => "00111111010111101000101100001010",
    211 => "01110001111110101100001011001111",
    212 => "01010111111010011110011110001001",
    213 => "00011111111011110000001101101100",
    214 => "01011110111101011110111011111000",
    215 => "01111010111010111001101111001011",
    216 => "01001111111111110100110110100010",
    217 => "01111111001111110011001111110111",
    218 => "01101110111111110111100111000001",
    219 => "01100111111101111001010101011001",
    220 => "01111110110011100110111010001110",
    221 => "00111111111111001010111100000011",
    222 => "01110110110010110101011000010110",
    223 => "01100111111011111000011010001010",
    224 => "01101101111111111011011000011110",
    225 => "00011111100111111101001100011011",
    226 => "00111010111011010100100100100011",
    227 => "01011110111111111101111011011110",
    228 => "01001101111111100101100101110011",
    229 => "00110111011101111101010101110100",
    230 => "01110011111111110111010110000011",
    231 => "01011111101111111000111101001111",
    232 => "01100111010101110100000100101100",
    233 => "01111110111111110010111001000100",
    234 => "01001111111111110001001001000101",
    235 => "00110000110101111010000011000011",
    236 => "01001111110111100010100001100000",
    237 => "01111111011101101001111111000011",
    238 => "01101111111011100101011010001000",
    239 => "00101111101111110101111110010111",
    240 => "01111010101100110110111110100111",
    241 => "01111011110010110010011110111100",
    242 => "01011111101110111110110101011000",
    243 => "01110110110110110000010101011010",
    244 => "01011010110111111101010001110001",
    245 => "01001011111101011100101100110010",
    246 => "01011010110111110100110000001110",
    247 => "01011101001111110000110100011010",
    248 => "00111011110111100001110111000111",
    249 => "00110001110111100100100000101001",
    250 => "01111000111111011111111011111100",
    251 => "01110111110111001011000011011111",
    252 => "01011010111000110011100010110011",
    253 => "00111111011110111010010111010010",
    254 => "01010101111011110111011011110001",
    255 => "01110111101110111001101111100001",
    256 => "01100111100111110011100000011101",
    257 => "00101101011101111001111101100011",
    258 => "00100110101111101100101000111000",
    259 => "00111110111110100110110001000000",
    260 => "01110111111101100111111110001101",
    261 => "01101011101110111110100010011111",
    262 => "01111101111110011001000111110011",
    263 => "00111111111111100101100011010110",
    264 => "00110010011101101101111111000110",
    265 => "01111101101101111000100111101100",
    266 => "01110110100111110101011101110000",
    267 => "01111111010101101110000101001000",
    268 => "01011000001111110101000111011010",
    269 => "01111101101111110000001010101100",
    270 => "01111111001101011011000101011000",
    271 => "01111011111110010110000000111110",
    272 => "01011110111111111000001011110011",
    273 => "01010010100100110001101000111011",
    274 => "01100011110110100000001111110000",
    275 => "01110111111100111100111000011100",
    276 => "00100110111111111111100010010011",
    277 => "01111111011100111100011111110010",
    278 => "01110111110111100101100110111111",
    279 => "01110001101011111011011000001001",
    280 => "01010111111100010001010001111101",
    281 => "01111111010111111010111001110010",
    282 => "01110001101111101110111110001011",
    283 => "00111110010111010101010000010010",
    284 => "00110101011010101110101111101000",
    285 => "01001101111111100000110010010010",
    286 => "01001111101011101000000011111011",
    287 => "01111011111101100001100010100101",
    288 => "00111100101101111001001000000110",
    289 => "01101010111110101001111000010000",
    290 => "00010110101011001011001001111001",
    291 => "01111011001111111000011100010101",
    292 => "01001111010101111100000001001111",
    293 => "01011110011111110001110101111010",
    294 => "01110111111001111010000011100101",
    295 => "00110101111101111100101100111110",
    296 => "01111010011111110001101110111001",
    297 => "01101111111010110010101011001111",
    298 => "01010111111101111000100010111100",
    299 => "00010111111011110111010100110101",
    300 => "01111110101110110110001011011101",
    301 => "01110111110110111001000101100111",
    302 => "01001111101111010001011011111110",
    303 => "00110110011110110100001010100111",
    304 => "01101111001001011110110100011010",
    305 => "01001111111111111010000001111010",
    306 => "01101011101111010011001110100100",
    307 => "01011111100110101110010101101001",
    308 => "01011001101111101111100011011000",
    309 => "00100011101101011100111011100101",
    310 => "01000110110111100010011011101111",
    311 => "00101111111111010001011011100100",
    312 => "00111011101111110011101001001011",
    313 => "01001111111100110000010101001111",
    314 => "01011111011011111111001010010100",
    315 => "00101001110100111111101100101011",
    316 => "01101111111011111110011111111000",
    317 => "00101111101100011010011110100101",
    318 => "01110111101111110100011110110010",
    319 => "01101100011011111000101011000001",
    320 => "01111110011001100010001010111110",
    321 => "01101110110111110101001111100110",
    322 => "00111001011011110101110011011111",
    323 => "01011101101101111100010100111001",
    324 => "01010100010111110100100110001000",
    325 => "01110010111101111101011101001100",
    326 => "01111110100111011111101001000100",
    327 => "01111100011111101101111000110111",
    328 => "01011101011010101001110011111011",
    329 => "00100111111101000010011000010000",
    330 => "01101101111101111001101010101001",
    331 => "01101011111111111010111110010100",
    332 => "01111010111111010110001001110101",
    333 => "00111101101101001100101010001001",
    334 => "01111110111011111111100010111011",
    335 => "01110111101111101110101101010011",
    336 => "00111000101111010101011110111110",
    337 => "01101001110011111010101101010010",
    338 => "00001111111111110100010010101011",
    339 => "01111100111111110001000110111110",
    340 => "00011100010010110111000011001111",
    341 => "00011110111111110010111101101001",
    342 => "01011111111010000000101110010110",
    343 => "01111100110110111011011100110110",
    344 => "01011111011011111110011100000011",
    345 => "01000111101011000010110110000110",
    346 => "01111101000111111010101011111101",
    347 => "01001101011110110110010000001000",
    348 => "00101111111100110001011101101111",
    349 => "00011011101011111001001010100110",
    350 => "01111101111111110100110100000000",
    351 => "00101101111111110110010111000101",
    352 => "00011111101101110010111010000111",
    353 => "01111011111100110100011000000101",
    354 => "01011111111101111001001110110110",
    355 => "00110100111011011001000000010111",
    356 => "00111111100001010110001111000110",
    357 => "01101111010111011001111100111101",
    358 => "01110111011111001100110100100000",
    359 => "00110110001000110001011111101110",
    360 => "01000111011111010011001110111011",
    361 => "00111101111111000010001010001110",
    362 => "00111011111111101110110000101010",
    363 => "00110111011010100100101000101001",
    364 => "01101111111011101111110011001011",
    365 => "00111111010100101011101000101001",
    366 => "00101110111011111100000100000110",
    367 => "00111110101111110101011111110010",
    368 => "00111111101110010101100101000001",
    369 => "01111010011111101110111000011011",
    370 => "00111111101111010010101100010101",
    371 => "01001011111110110100111011110010",
    372 => "00010110101011110110111101011111",
    373 => "01101101101011111000100001111000",
    374 => "00111111001101100110000101100101",
    375 => "01000111011110101110010100000100",
    376 => "01101111111011011100110001100001",
    377 => "01001001001111100001110011011100",
    378 => "01110111111101101101111100011100",
    379 => "01111101011011101111010001111110",
    380 => "00010011010100101101011100110101",
    381 => "01111111001111111111010011011110",
    382 => "01001110011111111100000110011110",
    383 => "00101111101110111110101011100000",
    384 => "00110111111111010100011010011101",
    385 => "00011111101100000110101011110101",
    386 => "01111010010101010101100011111000",
    387 => "01110111011101100001100000111101",
    388 => "01111101101110110111111110000100",
    389 => "00111110111011001000110001110111",
    390 => "01111001111111111100011100110011",
    391 => "00111111101101011100010111111110",
    392 => "01111010110110111010000010101001",
    393 => "01011101101111101011100111100001",
    394 => "00010111111101110001111111100111",
    395 => "00110111110101011110010001000000",
    396 => "00110111111111101100000000111101",
    397 => "00101011111111010110001011100100",
    398 => "01000110100011011100000100010010",
    399 => "00011111101010110011111100010001",
    400 => "01010111111011111001101011100010",
    401 => "01111010011111111111101101111011",
    402 => "00111111111111111101000011110010",
    403 => "00011101111111111101100011110011",
    404 => "00011110111111111111100101101110",
    405 => "00011011100111110010101110111001",
    406 => "00001011011111011000000111001101",
    407 => "01111011111011100001100111011100",
    408 => "01111011110110111101100110110111",
    409 => "01111101111111111100110011000100",
    410 => "01101101000101110100111010001000",
    411 => "00111011011111010110001111010110",
    412 => "01111001111111100011100000011111",
    413 => "01111011011111110101101011101101",
    414 => "00011110110111110001001100111100",
    415 => "00101110111111111111000101001110",
    416 => "01101110110010010010111101000101",
    417 => "00001111101111011001011010101010",
    418 => "00010101100110110101101001100101",
    419 => "00000110101111101010011100101010",
    420 => "00111010111111110010101000101111",
    421 => "01101101111011110000111010010111",
    422 => "01111010010011100110010010100101",
    423 => "01110001111011010111110111001110",
    424 => "01101111111111101010011001000101",
    425 => "01011111101110111011111001101011",
    426 => "01000010111110100111001010101111",
    427 => "01110111111111010101001001100011",
    428 => "01110101101110010001000110110000",
    429 => "00111111110110100010011000111101",
    430 => "01111100101101111000100111100000",
    431 => "00111101100011110011100001110011",
    432 => "01111110111111110000011011000000",
    433 => "00010101110111110101101000000010",
    434 => "00111101111111101111110110100101",
    435 => "01100011111111101111000000010001",
    436 => "01101110111111011111000011010011",
    437 => "01110111100011111010010100000110",
    438 => "00010100111111100100011101000101",
    439 => "01111101111101111010111100010100",
    440 => "01100101011111111001011110111010",
    441 => "00111001111010110001110111110001",
    442 => "01101111011111111000001100011111",
    443 => "01011111000011110101000111000100",
    444 => "01001110101101111100010011010000",
    445 => "01101011111100010011111000001011",
    446 => "01011100111111011110110011011010",
    447 => "00111111101111101110000011100111",
    448 => "01011110101111100101011010110101",
    449 => "01100110111011111011100000000100",
    450 => "00101100111111111000001001110111",
    451 => "01111101111111111111010101000011",
    452 => "01011111110010110001011101101101",
    453 => "01011111101110111010001000001100",
    454 => "01110001011101010010111100001100",
    455 => "01111110111101100001100010100111",
    456 => "00110110100111000101001010011000",
    457 => "01100011111101000111101011000111",
    458 => "00111010111100110100110000101100",
    459 => "01111101101011110000101100101000",
    460 => "01111110101111111011100011010000",
    461 => "00001111100001101100110010001110",
    462 => "01100101100110111100101010011100",
    463 => "01111101001100110101011001001101",
    464 => "01101111111110000010110101101010",
    465 => "01111101110101110111110110010000",
    466 => "01110100111111101010001110001001",
    467 => "01111101001111110111000010111101",
    468 => "01000111110101111101101110101100",
    469 => "01101011111111111111001011001001",
    470 => "01101101101101111001100100001110",
    471 => "01111011111111100000110111010001",
    472 => "01111011111111111010110100100111",
    473 => "01111101011011111001110010001001",
    474 => "01110101010111011001001100000011",
    475 => "01101110111110110110010011011111",
    476 => "01111011011011101110010000100011",
    477 => "00011011111111111011110000001110",
    478 => "00111111111111100000011010111101",
    479 => "01111100111101110101011001100100",
    480 => "01111001111111100101100100111010",
    481 => "01111101111110110000000101111110",
    482 => "01111101111110111011011000011110",
    483 => "01111110111001111000110101001110",
    484 => "00110110111111000010100100000111",
    485 => "01100111101111111010001000100010",
    486 => "01111110111011111001000011010101",
    487 => "00111111111111000111101111101110",
    488 => "01111101110111111001010000000100",
    489 => "01111011111101101000001101101001",
    490 => "01101111101111011000111101001000",
    491 => "01101011111101101011010000010000",
    492 => "01111110110111010111100100011010",
    493 => "01111111011111111000010011110100",
    494 => "01011111011111111010011101100101",
    495 => "00101110111110111100100101101100",
    496 => "01110101011111111000011000001101",
    497 => "00111111101111010010100001110010",
    498 => "01111101111111111110010111101100",
    499 => "01111110110000010000001010001001",
    500 => "01110111111110101001101010011001",
    501 => "01111110011111111100100110000110",
    502 => "01111101110111111000010110001111",
    503 => "01111110101110010111100101100100",
    504 => "01111110110110110011100001100100",
    505 => "00010111101101001101110010000111",
    506 => "00101101111011111000100010101100",
    507 => "00100111111110110111111001111011",
    508 => "00110101100001100001001111100111",
    509 => "01110001101111110001101001111100",
    510 => "00111101111101111111111101111100",
    511 => "01011110011100010010000100101000",
    512 => "01101111101011101101001100011000",
    513 => "01011101111001111100110001001110",
    514 => "01100111111111110110100001000101",
    515 => "01110100101010100101011101010000",
    516 => "01111101011110010100010000001011",
    517 => "01110011111110101000000001110011",
    518 => "01001001101001011011110100001100",
    519 => "01010110101010111010010101000001",
    520 => "01011111111111000001011111011010",
    521 => "01011101111111010001001110111100",
    522 => "01011110001111000111010101011001",
    523 => "00011011010011100111100101100011",
    524 => "01010111111001010001001100111100",
    525 => "01011111101111101101100111000110",
    526 => "01111110111111110100100011110110",
    527 => "01111100110111111011000011111001",
    528 => "01101101111011110111010010110110",
    529 => "01111101100001101100001011111010",
    530 => "00010111011001111110111010001100",
    531 => "01101111111111111111000101111110",
    532 => "00101110110011100010011110011000",
    533 => "01101110111110110111100000011111",
    534 => "01001111111111011000001010110101",
    535 => "00011110111100110010110000111101",
    536 => "00111001101101100110010110100010",
    537 => "01111111001001110010100010101010",
    538 => "00111011111011100010101011010111",
    539 => "00000101100111010111001011100101",
    540 => "00111011110111110100111010011111",
    541 => "01101111111011111101011111101010",
    542 => "01111100111001100111110011100000",
    543 => "01110011110101010001100010100110",
    544 => "01101110011111010100011011100000",
    545 => "01101111011111101001000010010101",
    546 => "01001000101111101011100010101111",
    547 => "00111011111001110011101101010001",
    548 => "01100111101111111001100010101110",
    549 => "01111110010100001101000111010111",
    550 => "01111010101011010000100100100101",
    551 => "01111011111111001101110101010101",
    552 => "01110011011110110011011001100111",
    553 => "00000101011001100011100010011001",
    554 => "01111100101111010000110000010110",
    555 => "01111110111110101000010010011111",
    556 => "01110111111111110001110101001100",
    557 => "01111110011101010011000010100000",
    558 => "01011001010011110100000101011010",
    559 => "01101000101110110111000111101011",
    560 => "00011011110101000101001101101100",
    561 => "00101100000111111111011010110011",
    562 => "00111011000111110000101100110100",
    563 => "01011111110111111001100110010100",
    564 => "00111110111111111010001000110010",
    565 => "01111110010001101101011010110110",
    566 => "01111111011011111100111111000011",
    567 => "01011011111101010100011101110100",
    568 => "01111101111011001011111111011010",
    569 => "01110010111110100101010101100101",
    570 => "01111110111111111011010100010101",
    571 => "01101111001111100011100111000001",
    572 => "01111101011011110001111011111010",
    573 => "00111111111011100010100110000000",
    574 => "01110100101101011001100101001001",
    575 => "01101100111110110100011110110011",
    576 => "01110111010111111101100010010111",
    577 => "01111010111111101111101000100001",
    578 => "01101111111111011000010000000000",
    579 => "01111010111111111111101001010010",
    580 => "01111111001111010101100000111001",
    581 => "01110111110110010111101101100101",
    582 => "01111000111010100001011000111010",
    583 => "01111011010011110101011001000011",
    584 => "01010010000001000110011110001010",
    585 => "00100110110011011111001001010000",
    586 => "01011111110100110001110100110010",
    587 => "01111110111110111001110000110010",
    588 => "01111011111001010101000010000101",
    589 => "01111111010111011001011101000100",
    590 => "01011111011111111100010100101100",
    591 => "01001011111011111010001111100111",
    592 => "01011110101111011001111101011111",
    593 => "01110111110111101010001111100011",
    594 => "01101101111011010110100001001110",
    595 => "01001111101111000001111100011000",
    596 => "01111010111111111011111101100011",
    597 => "01110101111111110111010000000101",
    598 => "01011111010111110110101101001000",
    599 => "01110110110101101010000011101101",
    600 => "01111111001111010101101001001100",
    601 => "01110111011111100101100101010111",
    602 => "01111101110011011010111100001101",
    603 => "01011101101111111101100101101111",
    604 => "01110110000101111110011111001000",
    605 => "01111011101111000110101011010000",
    606 => "01011111000111111110110110011011",
    607 => "00001100101101111001100110010101",
    608 => "01011010111110011110000101011010",
    609 => "01110111111111111010011100110001",
    610 => "01010110111111110010111010010110",
    611 => "01011111101100110001111110100111",
    612 => "01111011111101001110010101001100",
    613 => "00111110101011110110001011000000",
    614 => "00010011110011101111000101110010",
    615 => "00111111011011010011010000101101",
    616 => "00111101111111010001000101100001",
    617 => "00111111111111011110010010101010",
    618 => "00111011111011111010110000110111",
    619 => "00110101100011110000011010101000",
    620 => "00011110111011110001111110101100",
    621 => "01111001011001010100010010010110",
    622 => "01110111111110010010101110011110",
    623 => "01011010110110010001001000111010",
    624 => "01001100110110110111101101010000",
    625 => "01011111111111111110010101001010",
    626 => "01001110110111100001000001010100",
    627 => "01110111101101110001010011101011",
    628 => "01001111110111100000100100111010",
    629 => "01111101111101111000010011100011",
    630 => "00010110110011010010010111001010",
    631 => "00001111011101100100101100000011",
    632 => "01110111101111101101000001010101",
    633 => "01110111111111110100010111000001",
    634 => "01111010111011110100100001110101",
    635 => "00011101010011111001010111111100",
    636 => "01100001110111110110010000101000",
    637 => "01110111111111111011001011111011",
    638 => "01101110110111111001010001101011",
    639 => "01111011101111111011011100110011",
    640 => "01100111110011011100100101000011",
    641 => "01111110111011110100010001001011",
    642 => "01101111110101010011101010011101",
    643 => "01001010111111101000101011101100",
    644 => "01010111111011110101010111000100",
    645 => "00111110001110010001010011001010",
    646 => "01011010101111101100110100101010",
    647 => "01111111011001011111110100010110",
    648 => "01001111110010111101000110011101",
    649 => "01101111100111100000001101001011",
    650 => "01100111011101111101001010010110",
    651 => "01111101101111010010100100110101",
    652 => "01111101101001111101110111010101",
    653 => "00011101001111111011001111011101",
    654 => "01111101101000100011011101010101",
    655 => "01010111011011100101101101001110",
    656 => "01110110101100110101011010101110",
    657 => "01101100011110110100101000110001",
    658 => "01011110111111000010101000000010",
    659 => "01110111101111101101001010001011",
    660 => "00011111001001010100111110010000",
    661 => "01011011111111110001010100101100",
    662 => "01101111111001111111001010111111",
    663 => "00011011111111101011101001001110",
    664 => "00011010001111010110110101010011",
    665 => "01101001011111001101100110010100",
    666 => "01010001111011010010110100101101",
    667 => "00101001111111101001111001010000",
    668 => "01111011100111111000110010001010",
    669 => "01010101111101010010000011101100",
    670 => "00011111111010111010100111000010",
    671 => "01111110110111111110001010100111",
    672 => "01011100111111111100101011110000",
    673 => "01011011100011011100011000111000",
    674 => "01011011111111000010011101010101",
    675 => "01011010010101000110110101011100",
    676 => "01110111111110111100001100100110",
    677 => "01110100011111010011011000001001",
    678 => "01001111110111011011111111001111",
    679 => "01111110111111110101000110101010",
    680 => "00111111111100010111011010111010",
    681 => "00111111101001101110100110011001",
    682 => "00110111111100110000001011000001",
    683 => "00101111111011110000111101000000",
    684 => "00110011110111001010011010111111",
    685 => "01011101011011101000000001001000",
    686 => "01101011001110100010100111100011",
    687 => "01110000000110110010010110010110",
    688 => "01101100111111110110010110111001",
    689 => "01010111100101111100101101111111",
    690 => "00001110111011110110011011111111",
    691 => "00111101001011001111101011000001",
    692 => "00111011111110001011111100011110",
    693 => "00010100111111011010110010100110",
    694 => "01001111101011011010011110001100",
    695 => "01011111011101100000000011000011",
    696 => "01111111011111100111101000111110",
    697 => "01111110111111111011010111101100",
    698 => "01100101111011000000110101110000",
    699 => "00110101111011110010100110000010",
    700 => "00111101111110101111100001111000",
    701 => "00100110011111110011110110010101",
    702 => "01101111001111111111010100000011",
    703 => "01111110111111100001001001110110",
    704 => "01111101111111111011000000010110",
    705 => "00111111111101110010110111010010",
    706 => "00111111111100110110110010011010",
    707 => "01101011101111011011010000011110",
    708 => "01110011110101001110001100100011",
    709 => "00111011101011110011110010000001",
    710 => "00111111011011100010110111110001",
    711 => "00101101011011111010100011110101",
    712 => "01111110111010010010011110100000",
    713 => "01111101110100100010010100101110",
    714 => "01011110110001011110100100111111",
    715 => "00100111110101011111100001111011",
    716 => "01101101011111100011111011100000",
    717 => "00111110011111110100100000111011",
    718 => "01110110010111110010111101001011",
    719 => "00111011111101110101000100101101",
    720 => "01000101110010111001111010100001",
    721 => "01000011110011011100011110011110",
    722 => "00001111000111110110011000010000",
    723 => "00110110010100010000110001110100",
    724 => "01110111011011110100000101100011",
    725 => "01111001101111110011110000110001",
    726 => "01111111010111110001010001001011",
    727 => "00111101111111001001111000010100",
    728 => "00101111010111111011000000010000",
    729 => "00111000101111110101010011011110",
    730 => "00110111111111111010111000101000",
    731 => "01111101001011011001011000001010",
    732 => "01011111011111011110010100010101",
    733 => "00011100011001000111001001000000",
    734 => "01011111011011110101010001010011",
    735 => "01110111111111101100100010111000",
    736 => "00111110111011110111010010111000",
    737 => "01110011101011010111110000000011",
    738 => "00111111011101111100001011001010",
    739 => "01111110111111110011011010010110",
    740 => "01011110111001110010011001101001",
    741 => "01101101111111110110000001011010",
    742 => "01010100011010111000001100111001",
    743 => "01011000000101110100101111010001",
    744 => "01111101111110111011100011110111",
    745 => "01011111111110110110101111010110",
    746 => "01011011111110110011001000100010",
    747 => "01100110111110100010110101000111",
    748 => "01101111110111100110010101001011",
    749 => "01010101111100010110011111001111",
    750 => "01101101010111111000110101110101",
    751 => "00011101011111100101111101010000",
    752 => "00110110010110100110101001110011",
    753 => "00101011001011111100011011011110",
    754 => "01101101011011000010000100010101",
    755 => "01101101111100001110101111101010",
    756 => "01111101111111101001000111011011",
    757 => "01101110111100110100011100111011",
    758 => "00110011011111011111011110010000",
    759 => "01101011101110111001100111010011",
    760 => "01010111001111100000001111111100",
    761 => "01111111011011100111111011011001",
    762 => "01101101010111100110011001101100",
    763 => "01011111111111011010011010001001",
    764 => "01010000111111010001010111000111",
    765 => "00101000111111011011001000000101",
    766 => "00111111111011111100100111101101",
    767 => "01011100111110010000110100010010",
    768 => "01111101111011110111100101001001",
    769 => "01111101111110110110011100001010",
    770 => "01111011111111110000011101011110",
    771 => "01101011011110111001101010001100",
    772 => "01101101111001111100011111111000",
    773 => "00010111111011100111010010100010",
    774 => "01110111011110111001111010000101",
    775 => "01000110111110111100110111101111",
    776 => "01111111011110001111111111001001",
    777 => "01110111101101111100101010101111",
    778 => "00111010111111111000010101110100",
    779 => "00110111011110011111001000110110",
    780 => "01110111110110011101010101101000",
    781 => "01111011111111110011011111010110",
    782 => "00110011111010110110001000001000",
    783 => "01001111111111110011011011001000",
    784 => "00111110011011100010000111111001",
    785 => "00111101111011111100100111110000",
    786 => "00011101111010010100100110000001",
    787 => "01010011111111101010001010010100",
    788 => "01110000100110111011000110011110",
    789 => "00111011111111111110010011111011",
    790 => "01111111011111111100011011111000",
    791 => "01111101111011100100010111010011",
    792 => "01010011010011111010000111101000",
    793 => "01101101001010110100011100010111",
    794 => "00111011001111010101100111001011",
    795 => "00111110110110110101111001001000",
    796 => "01000010111101010111001000110010",
    797 => "00111101101111111100111010111001",
    798 => "01011011111110110011110011000111",
    799 => "01111101111111111100111000001010",
    800 => "01111000110111111101011001011101",
    801 => "01101110101111111110000100100010",
    802 => "01110111110111110011100101100011",
    803 => "00101101011111111000000110000100",
    804 => "01010111111110000011000010001101",
    805 => "01011011111101101011100110001001",
    806 => "01111110110111111100100010011111",
    807 => "00101111111101110100100111000110",
    808 => "00101011100111011101110000000010",
    809 => "00111111010011111011100011010110",
    810 => "00111011111111010011010000100100",
    811 => "00000011110111111011101010001100",
    812 => "01111111010111110110011100101011",
    813 => "00111101111101100001101100011000",
    814 => "01111011011111100101100101000000",
    815 => "00001110111101110111100101110001",
    816 => "00110010110111000110110100010001",
    817 => "01111101101110111011001100101111",
    818 => "01101100101110111011010111101110",
    819 => "01111110110011110101000000011001",
    820 => "01111111011111110011110101110001",
    821 => "01111001100101111011000111100000",
    822 => "01111100011011110111001000100011",
    823 => "01011001011011110111010001110011",
    824 => "01111101111111110000111010000100",
    825 => "00111100011111111000000100000010",
    826 => "01111110011111110011101111011001",
    827 => "01101101111111110011101101010001",
    828 => "01011101011001101010110101001000",
    829 => "01111100011101111001011110000001",
    830 => "01011101011011110000011000001001",
    831 => "01010110011000101100110100110000",
    832 => "01101110111000111100101111111100",
    833 => "01011111011111111111000000000010",
    834 => "01111101111111111110000001011000",
    835 => "01011011111110001010000101011001",
    836 => "01110011011111101001111100001000",
    837 => "01111011111111011111111010100100",
    838 => "01101010111111111110110011001011",
    839 => "01111011011011111010001100001000",
    840 => "01100101000110110001111101100011",
    841 => "01011011001111101010111110101001",
    842 => "01101110111111110001111001111101",
    843 => "01001111110001110000010000100111",
    844 => "01111011111110110010110000111101",
    845 => "00111101000110111100111110001100",
    846 => "01010010100110010000111101010011",
    847 => "00110011111011111110110100000001",
    848 => "00001101111110101101010011000001",
    849 => "01011011111111011100010000101001",
    850 => "00110101111101001001111110000110",
    851 => "01011111110111100011010111001001",
    852 => "01011101001011011010110001000011",
    853 => "01011011111111100110011010011000",
    854 => "00001101110111111011000001101000",
    855 => "00111111101111110100011011100110",
    856 => "01111011011101110101000011011011",
    857 => "01111101111111010101000000111000",
    858 => "01111011111100110011001110110001",
    859 => "01000011001111010111011010000101",
    860 => "01111001111111111110111001100011",
    861 => "01110010101011100011101111010111",
    862 => "01111011111111011100001101100100",
    863 => "01111011111111110010001110000000",
    864 => "01101111110000110001110111101011",
    865 => "01110100111101110100111001011001",
    866 => "01111010101101110000100110011001",
    867 => "01011110011101101011001101010001",
    868 => "00110011100111110010110011011101",
    869 => "01100011110111101101011110001100",
    870 => "01111110111101010011110011011010",
    871 => "00111011001111110110001111001100",
    872 => "00101110111110100010011011000110",
    873 => "01000111011000110010100011110100",
    874 => "01011111010101111101011001100101",
    875 => "00110110111111110011001000000010",
    876 => "01111101011001100100100111100011",
    877 => "01101101011011111110110110011010",
    878 => "00111110111111000011110100100110",
    879 => "01101000111101111001000000001001",
    880 => "01111101111011100011101110101101",
    881 => "01101111111111111101101101101101",
    882 => "00011000010010101111010000010110",
    883 => "01001111101100101111001010001001",
    884 => "01101111111100110110100011011001",
    885 => "01011111101101010001100110110011",
    886 => "01010010011110010101101010100000",
    887 => "00100011110111111111001100111101",
    888 => "01101111101001111000001001111101",
    889 => "00110100011111110101101011101011",
    890 => "00101100110111111101101111011111",
    891 => "01101101111111111010100111100101",
    892 => "00111111011111000001001000110001",
    893 => "01011111111110101101010100000000",
    894 => "01101101100010011101010101100100",
    895 => "01110001011111011011100000101110",
    896 => "01010111101110111111111010101100",
    897 => "01110110111110100000000000010000",
    898 => "01110011110111111001101111100110",
    899 => "00101110101111111011111001100101",
    900 => "01011010100111100010000111111100",
    901 => "01001101111010010001100010010010",
    902 => "00111111110011110000000000110001",
    903 => "01011011010111011000111001000011",
    904 => "01111110011011110100111110001110",
    905 => "01111111011100111111111111101011",
    906 => "01011111110111010011001110011101",
    907 => "01001111111111111001000111101011",
    908 => "01100111110111110110000101110101",
    909 => "01011101101110110110110110100110",
    910 => "01111110111100100111100001100000",
    911 => "01111110111100011010110100111111",
    912 => "01101001011101110101111100010101",
    913 => "01111111011110110110101100001010",
    914 => "00111111001001110100110111100100",
    915 => "00011111110011101111010110010010",
    916 => "00101111111111000000100110100100",
    917 => "01011111111101011110001111101001",
    918 => "01111010101011101010100100110011",
    919 => "01110100111111111101110001001111",
    920 => "00111111111011101111001000110100",
    921 => "01101100111111110111011011111011",
    922 => "01111111011101010001100010001001",
    923 => "00100111101110001110101101101110",
    924 => "01100111111011111111001000010011",
    925 => "00011111011100101111001010000010",
    926 => "01010011111101111101110001000000",
    927 => "01010111011110101110100001110111",
    928 => "01111111010110110110111100010001",
    929 => "01100111111011101101010001010001",
    930 => "01011101111111010101010110100011",
    931 => "00111001100011110111001011001000",
    932 => "01011111111111001110011111001011",
    933 => "01011110111111011010101110111001",
    934 => "00101011110010110001010010111101",
    935 => "00101110111110101011000110011011",
    936 => "00111000100111101001011111110101",
    937 => "01110101111111111000101100010001",
    938 => "01111110111001010000000100000110",
    939 => "01110111110110100011011010101110",
    940 => "01111110111111000111101011001000",
    941 => "01010111111010111011000100111111",
    942 => "00000111111010110100111001111110",
    943 => "01000011110111101011000000100000",
    944 => "01010111111010110100000001101111",
    945 => "01110110110000101110010010101001",
    946 => "00111110011111010111010000110001",
    947 => "00001100101101101111100011110010",
    948 => "01111100111010111011111011011011",
    949 => "01110111011100111111101010000011",
    950 => "01110111110101111011001011111011",
    951 => "01100101111011010001110010000100",
    952 => "01011111111111101000101101100001",
    953 => "01101111101110111100000001001100",
    954 => "01101011100011100111100001101110",
    955 => "00111001111111111001000011101011",
    956 => "01101110001111011010001101110010",
    957 => "01001110111110111010010100000110",
    958 => "00111101111111110110000000101101",
    959 => "01111111001111110001111001011111",
    960 => "01111101101110110010010101011101",
    961 => "01110011111010111101110100100011",
    962 => "01011111111011101001110100011100",
    963 => "01010111010111111101010101010101",
    964 => "00110111111110111001010101111111",
    965 => "01110111110110111000100100100101",
    966 => "01001111110111011100000100010101",
    967 => "01011100111111111100011101010111",
    968 => "00111111111001011101100111110000",
    969 => "01111011111111110010100000000010",
    970 => "01011111011111101111100010100011",
    971 => "01111101101110111101100100001001",
    972 => "01111001001101110101001110001111",
    973 => "01111101111011111011011011100001",
    974 => "01111110111111111001001001010110",
    975 => "01111111011111110100111100101001",
    976 => "01101110010011011011111001000001",
    977 => "01010111100101100100011100011111",
    978 => "01110101110111001000010101101111",
    979 => "01001111111101000010101101110011",
    980 => "01111100101010000010011110100111",
    981 => "01101110111111110001100011100000",
    982 => "01111111011101100010111011000100",
    983 => "01100111111001110101110110101100",
    984 => "00111111111101111111110001111010",
    985 => "01010000010111111100010100010001",
    986 => "01111011111110110110111111101100",
    987 => "01000010011000111100000111110111",
    988 => "00011001111010000101100000110010",
    989 => "01111111011110110111000110111011",
    990 => "00111111111111101111110101100101",
    991 => "00111101111001101010101000001001",
    992 => "00111111111110111010110001110011",
    993 => "01010111111111110000101110011110",
    994 => "01110111110101010011111000001100",
    995 => "01111110111111011100010001101110",
    996 => "01001101011111110010001001000100",
    997 => "00100111111010101111111001111000",
    998 => "01111011111110100111100001101111",
    999 => "01111101100110011101111000100000");

  component fabs is
    port (A : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          Q : out std_logic_vector (31 downto 0));
  end component fabs;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (3 downto 0) of std_logic_vector (31 downto 0);
  signal cc : std_logic_vector (31 downto 0) := (others => '0');  
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0'); 
  signal Q_buff : std_logic_vector (7 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
  signal i_isRunning : std_logic := 'U';
  signal i_result : std_logic := '1';
begin  -- architecture fabs_tb

  i_fabs : fabs port map (s_a,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk,Q_buff) is
    variable ss : character;
    variable count : integer := 1;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      s_a <= a_lut (addr);
      cc <= ans_lut (addr);
      ccc <= cc ;

      if i_isRunning = '1' then  -- rising clock edge
        if ccc = c and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 1 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;

  end process ram_loop;

end architecture;
