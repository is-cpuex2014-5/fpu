library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity fadd_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity fadd_tb;

architecture testbench of fadd_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);

  constant a_lut : lut := (
    0 => "00000000000000000000000000000000",
    1 => "00000000000000000000000000000000",
    2 => "00111111011100000110011101110100",
    3 => "00000000000000000000000000000000",
    4 => "00111110101011110001011011100111",
    5 => "00111111010111001110100011000100",
    6 => "00000000000000000000000000000000",
    7 => "00111110111111111101010001001100",
    8 => "00111111010000011001110010011110",
    9 => "00000000000000000000000000000000",
    10 => "00111111001001000011010011100111",
    11 => "00000000000000000000000000000000",
    12 => "00111111010000011001110010011110",
    13 => "00000000000000000000000000000000",
    14 => "00111111001001000011010011100111",
    15 => "00000000000000000000000000000000",
    16 => "00000000000000000000000000000000",
    17 => "01000000000100000000000000000000",
    18 => "00000000000000000000000000000000",
    19 => "00000000000000000000000000000000",
    20 => "00000000000000000000000000000000",
    21 => "00000000000000000000000000000000",
    22 => "00000000000000000000000000000000",
    23 => "00000000000000000000000000000000",
    24 => "10111111000000100111001000100111",
    25 => "10111110000001011010100011000011",
    26 => "00000000000000000000000000000000",
    27 => "00111111011111011100111010000110",
    28 => "00111010111000110010111001111001",
    29 => "00000000000000000000000000000000",
    30 => "10111111000000100101110100000000",
    31 => "00111111011010110101000100110010",
    32 => "00000000000000000000000000000000",
    33 => "00111110110010000100010011011011",
    34 => "00111111000100000001101000110100",
    35 => "10111110001101001100110110101100",
    36 => "10111101101110011011111111100001",
    37 => "00000000000000000000000000000000",
    38 => "00111111011111101111000110110100",
    39 => "00111011101101000010101101100010",
    40 => "00000000000000000000000000000000",
    41 => "10111111000000100000010111110000",
    42 => "00111111011010010111011100101011",
    43 => "00000000000000000000000000000000",
    44 => "00111110110100001000011000001011",
    45 => "00111111000001111011101010011011",
    46 => "10111110001111000001011110011100",
    47 => "10111101101111001011111011001010",
    48 => "00000000000000000000000000000000",
    49 => "00111111011111101110100011100100",
    50 => "00111011101100001110010110000000",
    51 => "00000000000000000000000000000000",
    52 => "10111111000000100000100011101000",
    53 => "00111111011010011000001011100010",
    54 => "00000000000000000000000000000000",
    55 => "00111110110100000101001100011000",
    56 => "00111111000001111110100101011110",
    57 => "10111110001110111110110100110111",
    58 => "10111101101111001010110110111010",
    59 => "00000000000000000000000000000000",
    60 => "00111111011111101110100100010110",
    61 => "00111011101100001111100010000100",
    62 => "00000000000000000000000000000000",
    63 => "10111111000000100000100011010101",
    64 => "00111111011010011000001010100000",
    65 => "00000000000000000000000000000000",
    66 => "00111110110100000101010000111000",
    67 => "00111111000001111110100001010111",
    68 => "10111110001110111110111000100110",
    69 => "10111101101111001010111000011100",
    70 => "00000000000000000000000000000000",
    71 => "00111111011111101110100100010101",
    72 => "00111011101100001111100000011010",
    73 => "00000000000000000000000000000000",
    74 => "10111111000000100000100011010110",
    75 => "00111111011010011000001010100000",
    76 => "00000000000000000000000000000000",
    77 => "00111110110100000101010000110101",
    78 => "00111011101100001111100000011010",
    79 => "00111111000010010100101001000111",
    80 => "00000000000000000000000000000000",
    81 => "00000000000000000000000000000000",
    82 => "00000000000000000000000000000000",
    83 => "00000000000000000000000000000000",
    84 => "10111111000000100111001000100111",
    85 => "00111111011011000100001011110000",
    86 => "00000000000000000000000000000000",
    87 => "00111110110000111110010000011010",
    88 => "00111111000101010011011010101001",
    89 => "00000000000000000000000000000000",
    90 => "10111110001100001010010000100000",
    91 => "00111111001101011101010101100001",
    92 => "00000000000000000000000000000000",
    93 => "00111111001100000000110001110110",
    94 => "00111111010000001001011001100010",
    95 => "10111110000101000001011000101110",
    96 => "00111111001011100001010010111110",
    97 => "00000000000000000000000000000000",
    98 => "00111111001101111110101001010110",
    99 => "00111111001111011011000110010011",
    100 => "00000000000000000000000000000000",
    101 => "10111110000101011010111100100000",
    102 => "00111111001011101011110101000000",
    103 => "00000000000000000000000000000000",
    104 => "00111111001101110011100110010000",
    105 => "00111111001111011110001101000010",
    106 => "10111110000101011001001101101011",
    107 => "00111111001011101011000111100111",
    108 => "00000000000000000000000000000000",
    109 => "00111111001101110100010110000100",
    110 => "00111111001111011101111111111000",
    111 => "00000000000000000000000000000000",
    112 => "10111110000101011001010100111111",
    113 => "00111111001011101011001010101000",
    114 => "00000000000000000000000000000000",
    115 => "00111111001101110100010010111000",
    116 => "00111111001111011110000000110011",
    117 => "10111110000101011001010100100000",
    118 => "00111111001011101011001010011010",
    119 => "00000000000000000000000000000000",
    120 => "00111111001101110100010011000110",
    121 => "00111111001111011110000000101101",
    122 => "00000000000000000000000000000000",
    123 => "10111110000101011001010100100100",
    124 => "00111111001011101011001010011101",
    125 => "00000000000000000000000000000000",
    126 => "00111111001101110100010011000100",
    127 => "00111111001111011110000000110011",
    128 => "10111110000101011001010100100000",
    129 => "00111111001011101011001010011010",
    130 => "00000000000000000000000000000000",
    131 => "00111111001101110100010011000110",
    132 => "00111111001111011110000000101101",
    133 => "00000000000000000000000000000000",
    134 => "10111110000101011001010100100100",
    135 => "00111111001011101011001010011101",
    136 => "00000000000000000000000000000000",
    137 => "00111111001101110100010011000100",
    138 => "00111111001111011110000000101101",
    139 => "00111111101111011110000000110000",
    140 => "00000000000000000000000000000000",
    141 => "00000000000000000000000000000000",
    142 => "00000000000000000000000000000000",
    143 => "00000000000000000000000000000000",
    144 => "00000000000000000000000000000000",
    145 => "00000000000000000000000000000000",
    146 => "00000000000000000000000000000000",
    147 => "10111111000000100111001000100111",
    148 => "10111110110000111110010100101100",
    149 => "00000000000000000000000000000000",
    150 => "00111111011011000100001010110101",
    151 => "00111100100011001000110111100000",
    152 => "00000000000000000000000000000000",
    153 => "10111110111111111110001011001010",
    154 => "00111111011001010010111111000100",
    155 => "00000000000000000000000000000000",
    156 => "00111110111000100010011111010101",
    157 => "00111110111101110011101000110100",
    158 => "10111110010001111101000100010110",
    159 => "10111110100011110011111010111101",
    160 => "00000000000000000000000000000000",
    161 => "00111111011101011011010011110010",
    162 => "00111101010010101100010001110001",
    163 => "00000000000000000000000000000000",
    164 => "10111110111011010011111101001100",
    165 => "00111111010111111011011000101100",
    166 => "00000000000000000000000000000000",
    167 => "00111110111101100101011011111001",
    168 => "00111110111111011100001001010001",
    169 => "10111110010001001000000110011000",
    170 => "10111110100011100101011010001111",
    171 => "00000000000000000000000000000000",
    172 => "00111111011101011101011100100000",
    173 => "00111101010011000101111010111110",
    174 => "00000000000000000000000000000000",
    175 => "10111110111011010000000000011011",
    176 => "00111111010111111010110010001010",
    177 => "00000000000000000000000000000000",
    178 => "00111110111101100111100001111110",
    179 => "00111110111111100001001000100101",
    180 => "10111110010001000101100111011111",
    181 => "10111110100011100100101110010000",
    182 => "00000000000000000000000000000000",
    183 => "00111111011101011101100010111101",
    184 => "00111101010011000111000111111111",
    185 => "00000000000000000000000000000000",
    186 => "10111110111011001111110100100010",
    187 => "00111111010111111010110000010110",
    188 => "00000000000000000000000000000000",
    189 => "00111110111101100111101000010000",
    190 => "00111110111111100001010111100110",
    191 => "10111110010001000101100000000011",
    192 => "10111110100011100100101100001101",
    193 => "00000000000000000000000000000000",
    194 => "00111111011101011101100011010000",
    195 => "00111101010011000111001011101000",
    196 => "00000000000000000000000000000000",
    197 => "10111110111011001111110100000001",
    198 => "00111111010111111010110000010001",
    199 => "00000000000000000000000000000000",
    200 => "00111110111101100111101000100001",
    201 => "00111101010011000111001011101000",
    202 => "00111111000010111101001000111000",
    203 => "00000000000000000000000000000000",
    204 => "00000000000000000000000000000000",
    205 => "00111111000110011001100110011010",
    206 => "00000000000000000000000000000000",
    207 => "00000000000000000000000000000000",
    208 => "10111111000000100111001000100111",
    209 => "00111111010010010010101101110110",
    210 => "00000000000000000000000000000000",
    211 => "00111111000110111001011010010100",
    212 => "00111110001011011110101101111011",
    213 => "00000000000000000000000000000000",
    214 => "10111110101011010001001010010101",
    215 => "00111111010101111001110010010010",
    216 => "00000000000000000000000000000000",
    217 => "00111111000010000011110100110011",
    218 => "00111111001011100110011111110110",
    219 => "10111110000111101100011000110111",
    220 => "00111111000100001100010010000110",
    221 => "00000000000000000000000000000000",
    222 => "00111111010100011010001101111101",
    223 => "00111110101111001011001010000011",
    224 => "00000000000000000000000000000000",
    225 => "10111110011010111100000100001010",
    226 => "00111111010001110010001001000111",
    227 => "00000000000000000000000000000000",
    228 => "00111111000111011111111110000010",
    229 => "00111111010000011101100011000001",
    230 => "10111110000100110110011100011101",
    231 => "00111111000011001010111001111000",
    232 => "00000000000000000000000000000000",
    233 => "00111111010101001001001010011100",
    234 => "00111110101111100110111101101101",
    235 => "00000000000000000000000000000000",
    236 => "10111110011010100111110110111010",
    237 => "00111111010001101101100001010010",
    238 => "00000000000000000000000000000000",
    239 => "00111111000111100101010110100101",
    240 => "00111111010000011110010111000010",
    241 => "10111110000100110110000000010010",
    242 => "00111111000011001010101111010101",
    243 => "00000000000000000000000000000000",
    244 => "00111111010101001001010001110110",
    245 => "00111110101111100111000001100101",
    246 => "00000000000000000000000000000000",
    247 => "10111110011010100111110100000100",
    248 => "00111111010001101101100000101011",
    249 => "00000000000000000000000000000000",
    250 => "00111111000111100101010111010011",
    251 => "00111111010000011110010111010010",
    252 => "10111110000100110110000000001100",
    253 => "00111111000011001010101111010011",
    254 => "00000000000000000000000000000000",
    255 => "00111111010101001001010001111000",
    256 => "00111110101111100111000001110010",
    257 => "00000000000000000000000000000000",
    258 => "10111110011010100111110011111001",
    259 => "00111111010001101101100000101000",
    260 => "00000000000000000000000000000000",
    261 => "00111111000111100101010111010110",
    262 => "00111110101111100111000001110010",
    263 => "00111111100100001000111100000011",
    264 => "00000000000000000000000000000000",
    265 => "00000000000000000000000000000000",
    266 => "00000000000000000000000000000000",
    267 => "00000000000000000000000000000000",
    268 => "10111111000000100111001000100111",
    269 => "10111111000110111001011100001010",
    270 => "00000000000000000000000000000000",
    271 => "00111111010010010010101100010100",
    272 => "00111101011100010010110000001100",
    273 => "00000000000000000000000000000000",
    274 => "10111110111001110101001110001000",
    275 => "00111111010111101110010101110010",
    276 => "00000000000000000000000000000000",
    277 => "00111110111110010010011101111011",
    278 => "00111111000000101110001001011111",
    279 => "10111110010000001001101000001010",
    280 => "10111110111001011110001011111100",
    281 => "00000000000000000000000000000000",
    282 => "00111111011001000011100011101011",
    283 => "00111110000111100011011000100100",
    284 => "00000000000000000000000000000000",
    285 => "10111110101100111001000010110110",
    286 => "00111111010110001011011110101100",
    287 => "00000000000000000000000000000000",
    288 => "00111111000001101001000010101110",
    289 => "00111111001010100100001101000010",
    290 => "10111110001000010111000111100011",
    291 => "10111110110101101100001101100111",
    292 => "00000000000000000000000000000000",
    293 => "00111111011010000000000010101100",
    294 => "00111110001001110110011000111101",
    295 => "00000000000000000000000000000000",
    296 => "10111110101011111011011001110000",
    297 => "00111111010110000001001110010000",
    298 => "00000000000000000000000000000000",
    299 => "00111111000001111000101000010100",
    300 => "00111111001011001100001011011100",
    301 => "10111110000111111101001010111100",
    302 => "10111110110101011110001110011011",
    303 => "00000000000000000000000000000000",
    304 => "00111111011010000011010111111111",
    305 => "00111110001001111101110100011111",
    306 => "00000000000000000000000000000000",
    307 => "10111110101011111000010110100101",
    308 => "00111111010110000000101100101000",
    309 => "00000000000000000000000000000000",
    310 => "00111111000001111001011011000111",
    311 => "00111111001011001110000111001000",
    312 => "10111110000111111011111011011101",
    313 => "10111110110101011101100011010101",
    314 => "00000000000000000000000000000000",
    315 => "00111111011010000011100010001110",
    316 => "00111110001001111110001011000101",
    317 => "00000000000000000000000000000000",
    318 => "10111110101011111000001101010100",
    319 => "00111111010110000000101011000010",
    320 => "00000000000000000000000000000000",
    321 => "00111111000001111001011101100000",
    322 => "00111110001001111110001011000101",
    323 => "00111111010101101101101111110011",
    324 => "00000000000000000000000000000000",
    325 => "00000000000000000000000000000000",
    326 => "00111110110011001100110011001110",
    327 => "00000000000000000000000000000000",
    328 => "00000000000000000000000000000000",
    329 => "10111111000000100111001000100111",
    330 => "00111111000110111001011100001100",
    331 => "00000000000000000000000000000000",
    332 => "00111111010010010010101100010010",
    333 => "00111101011100010010110000011000",
    334 => "00000000000000000000000000000000",
    335 => "10111110111001110101001110001000",
    336 => "00111111010111101110010101110010",
    337 => "00000000000000000000000000000000",
    338 => "00111110111110010010011101111011",
    339 => "00111111000000101110001001100000",
    340 => "10111110010000001001101000001010",
    341 => "00111110111001011110001011111111",
    342 => "00000000000000000000000000000000",
    343 => "00111111011001000011100011101010",
    344 => "00111110000111100011011000101100",
    345 => "00000000000000000000000000000000",
    346 => "10111110101100111001000010110011",
    347 => "00111111010110001011011110101011",
    348 => "00000000000000000000000000000000",
    349 => "00111111000001101001000010110000",
    350 => "00111111001010100100001101000010",
    351 => "10111110001000010111000111100011",
    352 => "00111110110101101100001101101010",
    353 => "00000000000000000000000000000000",
    354 => "00111111011010000000000010101100",
    355 => "00111110001001110110011001000000",
    356 => "00000000000000000000000000000000",
    357 => "10111110101011111011011001101100",
    358 => "00111111010110000001001110010001",
    359 => "00000000000000000000000000000000",
    360 => "00111111000001111000101000010010",
    361 => "00111111001011001100001011100100",
    362 => "10111110000111111101001010111001",
    363 => "00111110110101011110001110011100",
    364 => "00000000000000000000000000000000",
    365 => "00111111011010000011010111111110",
    366 => "00111110001001111101110100101011",
    367 => "00000000000000000000000000000000",
    368 => "10111110101011111000010110100001",
    369 => "00111111010110000000101100100111",
    370 => "00000000000000000000000000000000",
    371 => "00111111000001111001011011001000",
    372 => "00111111001011001110000111001010",
    373 => "10111110000111111011111011011101",
    374 => "00111110110101011101100011011000",
    375 => "00000000000000000000000000000000",
    376 => "00111111011010000011100010001101",
    377 => "00111110001001111110001011001100",
    378 => "00000000000000000000000000000000",
    379 => "10111110101011111000001101001111",
    380 => "00111111010110000000101011000010",
    381 => "00000000000000000000000000000000",
    382 => "00111111000001111001011101100000",
    383 => "00111110001001111110001011001100",
    384 => "00111111010101101101101111111010",
    385 => "00000000000000000000000000000000",
    386 => "00000000000000000000000000000000",
    387 => "00000000000000000000000000000000",
    388 => "00000000000000000000000000000000",
    389 => "00000000000000000000000000000000",
    390 => "00000000000000000000000000000000",
    391 => "00000000000000000000000000000000",
    392 => "10111111000000100111001000100111",
    393 => "10111111010010011011111110010110",
    394 => "00000000000000000000000000000000",
    395 => "00111111000101001000011110100000",
    396 => "00111110001011011110101111000010",
    397 => "00000000000000000000000000000000",
    398 => "10111110101011010001001001111000",
    399 => "00111111010101111001110010001110",
    400 => "00000000000000000000000000000000",
    401 => "00111111000010000011110100111010",
    402 => "00111111001011100110100000001010",
    403 => "10111110000111101100011000101000",
    404 => "10111111000100001100010010000010",
    405 => "00000000000000000000000000000000",
    406 => "00111111010100011010001110000000",
    407 => "00111110101111001011001010001010",
    408 => "00000000000000000000000000000000",
    409 => "10111110011010111100000100000101",
    410 => "00111111010001110010001001000110",
    411 => "00000000000000000000000000000000",
    412 => "00111111000111011111111110000011",
    413 => "00111111010000011101100011000001",
    414 => "10111110000100110110011100011101",
    415 => "10111111000011001010111001110111",
    416 => "00000000000000000000000000000000",
    417 => "00111111010101001001001010011110",
    418 => "00111110101111100110111101100011",
    419 => "00000000000000000000000000000000",
    420 => "10111110011010100111110110111111",
    421 => "00111111010001101101100001010101",
    422 => "00000000000000000000000000000000",
    423 => "00111111000111100101010110100010",
    424 => "00111111010000011110010111001001",
    425 => "10111110000100110110000000010010",
    426 => "10111111000011001010101111010100",
    427 => "00000000000000000000000000000000",
    428 => "00111111010101001001010001110111",
    429 => "00111110101111100111000001101010",
    430 => "00000000000000000000000000000000",
    431 => "10111110011010100111110100000010",
    432 => "00111111010001101101100000101000",
    433 => "00000000000000000000000000000000",
    434 => "00111111000111100101010111010110",
    435 => "00111111010000011110010111001000",
    436 => "10111110000100110110000000010010",
    437 => "10111111000011001010101111010100",
    438 => "00000000000000000000000000000000",
    439 => "00111111010101001001010001110111",
    440 => "00111110101111100111000001101010",
    441 => "00000000000000000000000000000000",
    442 => "10111110011010100111110100000010",
    443 => "00111111010001101101100000101000",
    444 => "00000000000000000000000000000000",
    445 => "00111111000111100101010111010110",
    446 => "00111110101111100111000001101010",
    447 => "00111111100100001000111011111110",
    448 => "00000000000000000000000000000000",
    449 => "00000000000000000000000000000000",
    450 => "00111110010011001100110011001110",
    451 => "00000000000000000000000000000000",
    452 => "00000000000000000000000000000000",
    453 => "10111111000000100111001000100111",
    454 => "00111110110000111110010100101110",
    455 => "00000000000000000000000000000000",
    456 => "00111111011011000100001010110101",
    457 => "00111100100011001000110111100010",
    458 => "00000000000000000000000000000000",
    459 => "10111110111111111110001011001010",
    460 => "00111111011001010010111111000100",
    461 => "00000000000000000000000000000000",
    462 => "00111110111000100010011111010101",
    463 => "00111110111101110011101000110111",
    464 => "10111110010001111101000100010110",
    465 => "00111110100011110011111010111111",
    466 => "00000000000000000000000000000000",
    467 => "00111111011101011011010011110010",
    468 => "00111101010010101100010001111000",
    469 => "00000000000000000000000000000000",
    470 => "10111110111011010011111101001001",
    471 => "00111111010111111011011000101100",
    472 => "00000000000000000000000000000000",
    473 => "00111110111101100101011011111001",
    474 => "00111110111111011100001001010011",
    475 => "10111110010001001000000110011000",
    476 => "00111110100011100101011010010001",
    477 => "00000000000000000000000000000000",
    478 => "00111111011101011101011100100000",
    479 => "00111101010011000101111011000101",
    480 => "00000000000000000000000000000000",
    481 => "10111110111011010000000000011000",
    482 => "00111111010111111010110010001010",
    483 => "00000000000000000000000000000000",
    484 => "00111110111101100111100001111110",
    485 => "00111110111111100001001000101000",
    486 => "10111110010001000101100111011111",
    487 => "00111110100011100100101110010010",
    488 => "00000000000000000000000000000000",
    489 => "00111111011101011101100010111101",
    490 => "00111101010011000111001000001000",
    491 => "00000000000000000000000000000000",
    492 => "10111110111011001111110100100010",
    493 => "00111111010111111010110000010110",
    494 => "00000000000000000000000000000000",
    495 => "00111110111101100111101000010000",
    496 => "00111110111111100001010111101001",
    497 => "10111110010001000101100000000011",
    498 => "00111110100011100100101100001111",
    499 => "00000000000000000000000000000000",
    500 => "00111111011101011101100011010000",
    501 => "00111101010011000111001011101111",
    502 => "00000000000000000000000000000000",
    503 => "10111110111011001111110011111110",
    504 => "00111111010111111010110000010000",
    505 => "00000000000000000000000000000000",
    506 => "00111110111101100111101000100100",
    507 => "00111101010011000111001011101111",
    508 => "00111111000010111101001000111011",
    509 => "00000000000000000000000000000000",
    510 => "00000000000000000000000000000000",
    511 => "00000000000000000000000000000000",
    512 => "00000000000000000000000000000000",
    513 => "10111111000000100111001000100111",
    514 => "10111111011001111101010001000010",
    515 => "00000000000000000000000000000000",
    516 => "00111110100111001011000010111000",
    517 => "00111111000101010011111100101100",
    518 => "00000000000000000000000000000000",
    519 => "10111110001100001001110101011111",
    520 => "00111111001101011101001011100010",
    521 => "00000000000000000000000000000000",
    522 => "00111111001100000000111011001011",
    523 => "00111111010000001001010111011100",
    524 => "10111110000101000001011001110110",
    525 => "10111111001011100001010011011100",
    526 => "00000000000000000000000000000000",
    527 => "00111111001101111110101000110110",
    528 => "00111111001111011011000110010111",
    529 => "00000000000000000000000000000000",
    530 => "10111110000101011010111100011110",
    531 => "00111111001011101011110100111111",
    532 => "00000000000000000000000000000000",
    533 => "00111111001101110011100110010010",
    534 => "00111111001111011110001100111111",
    535 => "10111110000101011001001101101011",
    536 => "10111111001011101011000111100111",
    537 => "00000000000000000000000000000000",
    538 => "00111111001101110100010110000100",
    539 => "00111111001111011101111111110101",
    540 => "00000000000000000000000000000000",
    541 => "10111110000101011001010101000011",
    542 => "00111111001011101011001010101010",
    543 => "00000000000000000000000000000000",
    544 => "00111111001101110100010010110110",
    545 => "00111111001111011110000000111010",
    546 => "10111110000101011001010100011010",
    547 => "10111111001011101011001010010110",
    548 => "00000000000000000000000000000000",
    549 => "00111111001101110100010011001011",
    550 => "00111111001111011110000000100011",
    551 => "00000000000000000000000000000000",
    552 => "10111110000101011001010100100111",
    553 => "00111111001011101011001010011110",
    554 => "00000000000000000000000000000000",
    555 => "00111111001101110100010011000011",
    556 => "00111111001111011110000000101101",
    557 => "10111110000101011001010100100100",
    558 => "10111111001011101011001010011011",
    559 => "00000000000000000000000000000000",
    560 => "00111111001101110100010011000110",
    561 => "00111111001111011110000000101010",
    562 => "00000000000000000000000000000000",
    563 => "10111110000101011001010100100100",
    564 => "00111111001011101011001010011101",
    565 => "00000000000000000000000000000000",
    566 => "00111111001101110100010011000100",
    567 => "00111111001111011110000000101010",
    568 => "00111111101111011110000000101110",
    569 => "00000000000000000000000000000000",
    570 => "00000000000000000000000000000000",
    571 => "00000000000000000000000000000000",
    572 => "00000000000000000000000000000000",
    573 => "00000000000000000000000000000000",
    574 => "10111111000000100111001000100111",
    575 => "00111110000001011010100011000011",
    576 => "00000000000000000000000000000000",
    577 => "00111111011111011100111010000110",
    578 => "00111010111000110010111001111001",
    579 => "00000000000000000000000000000000",
    580 => "10111111000000100101110100000000",
    581 => "00111111011010110101000100110010",
    582 => "00000000000000000000000000000000",
    583 => "00111110110010000100010011011011",
    584 => "00111111000100000001101000110100",
    585 => "10111110001101001100110110101100",
    586 => "00111101101110011011111111100001",
    587 => "00000000000000000000000000000000",
    588 => "00111111011111101111000110110100",
    589 => "00111011101101000010101101100010",
    590 => "00000000000000000000000000000000",
    591 => "10111111000000100000010111110000",
    592 => "00111111011010010111011100101011",
    593 => "00000000000000000000000000000000",
    594 => "00111110110100001000011000001011",
    595 => "00111111000001111011101010011011",
    596 => "10111110001111000001011110011100",
    597 => "00111101101111001011111011001010",
    598 => "00000000000000000000000000000000",
    599 => "00111111011111101110100011100100",
    600 => "00111011101100001110010110000000",
    601 => "00000000000000000000000000000000",
    602 => "10111111000000100000100011101000",
    603 => "00111111011010011000001011100010",
    604 => "00000000000000000000000000000000",
    605 => "00111110110100000101001100011000",
    606 => "00111111000001111110100101011110",
    607 => "10111110001110111110110100110111",
    608 => "00111101101111001010110110111010",
    609 => "00000000000000000000000000000000",
    610 => "00111111011111101110100100010110",
    611 => "00111011101100001111100010000100",
    612 => "00000000000000000000000000000000",
    613 => "10111111000000100000100011010101",
    614 => "00111111011010011000001010100000",
    615 => "00000000000000000000000000000000",
    616 => "00111110110100000101010000111000",
    617 => "00111111000001111110100001010111",
    618 => "10111110001110111110111000100110",
    619 => "00111101101111001010111000011100",
    620 => "00000000000000000000000000000000",
    621 => "00111111011111101110100100010101",
    622 => "00111011101100001111100000011010",
    623 => "00000000000000000000000000000000",
    624 => "10111111000000100000100011010110",
    625 => "00111111011010011000001010100000",
    626 => "00000000000000000000000000000000",
    627 => "00111110110100000101010000110101",
    628 => "00111011101100001111100000011010",
    629 => "00111111000010010100101001000111",
    630 => "00000000000000000000000000000000",
    631 => "00000000000000000000000000000000",
    632 => "00000000000000000000000000000000",
    633 => "00000000000000000000000000000000",
    634 => "00000000000000000000000000000000",
    635 => "00000000000000000000000000000000",
    636 => "00000000000000000000000000000000",
    637 => "10111111000000100111001000100111",
    638 => "10111110000001011010100010111011",
    639 => "00000000000000000000000000000000",
    640 => "00111111011111011100111010000110",
    641 => "00111010111000110010111001011111",
    642 => "00000000000000000000000000000000",
    643 => "10111111000000100101110100000000",
    644 => "00111111010001111111010000001011",
    645 => "00000000000000000000000000000000",
    646 => "00111111000111010000100101010000",
    647 => "00111110001010111011101101011010",
    648 => "10111110101011011111001100101101",
    649 => "10111101111001010110001010101010",
    650 => "00000000000000000000000000000000",
    651 => "00111111011111100110001100110010",
    652 => "00111011010111101110010001111000",
    653 => "00000000000000000000000000000000",
    654 => "10111111000000100011110011110011",
    655 => "00111111010001101101110111110101",
    656 => "00000000000000000000000000000000",
    657 => "00111111000111100100111100011000",
    658 => "00111110001010100000010011001011",
    659 => "10111110101011101010010010010100",
    660 => "10111101111001011001001111111110",
    661 => "00000000000000000000000000000000",
    662 => "00111111011111100110001001111111",
    663 => "00111011010111011110000001100111",
    664 => "00000000000000000000000000000000",
    665 => "10111111000000100011110101001011",
    666 => "00111111010001101110000001110100",
    667 => "00000000000000000000000000000000",
    668 => "00111111000111100100110000110001",
    669 => "00111110001010100000100001110111",
    670 => "10111110101011101010001100010011",
    671 => "10111101111001011001001110010101",
    672 => "00000000000000000000000000000000",
    673 => "00111111011111100110001010000000",
    674 => "00111011010111011110001010011010",
    675 => "00000000000000000000000000000000",
    676 => "10111111000000100011110101001010",
    677 => "00111111010001101110000001101111",
    678 => "00000000000000000000000000000000",
    679 => "00111111000111100100110000110111",
    680 => "00111110001010100000100001110010",
    681 => "10111110101011101010001100011000",
    682 => "10111101111001011001001110010101",
    683 => "00000000000000000000000000000000",
    684 => "00111111011111100110001010000000",
    685 => "00111011010111011110001010010010",
    686 => "00000000000000000000000000000000",
    687 => "10111111000000100011110101001010",
    688 => "00111111010001101110000001101111",
    689 => "00000000000000000000000000000000",
    690 => "00111111000111100100110000110111",
    691 => "00111011010111011110001010010010",
    692 => "00111110001011010111111111111100",
    693 => "00000000000000000000000000000000",
    694 => "00000000000000000000000000000000",
    695 => "00111111010011001100110011001110",
    696 => "00000000000000000000000000000000",
    697 => "00000000000000000000000000000000",
    698 => "10111111000000100111001000100111",
    699 => "00111111011011000100001011110000",
    700 => "00000000000000000000000000000000",
    701 => "00111110110000111110010000010110",
    702 => "00111111000101010011011010101111",
    703 => "00000000000000000000000000000000",
    704 => "10111110001100001010010000011001",
    705 => "00111111000101101000101111111010",
    706 => "00000000000000000000000000000000",
    707 => "00111111010011010011111101011011",
    708 => "00111110101110011001111010001110",
    709 => "10111110011011100000011010100101",
    710 => "00111111010001111010010101101000",
    711 => "00000000000000000000000000000000",
    712 => "00111111000111010110010111101111",
    713 => "00111111010000011011111011011111",
    714 => "00000000000000000000000000000000",
    715 => "10111110000100110111010100011000",
    716 => "00111111000011001011001110110100",
    717 => "00000000000000000000000000000000",
    718 => "00111111010101001000111011110000",
    719 => "00111110101111100110110101011010",
    720 => "10111110011010100111111100111000",
    721 => "00111111010001101101100010101100",
    722 => "00000000000000000000000000000000",
    723 => "00111111000111100101010100111101",
    724 => "00111111010000011110010110111101",
    725 => "00000000000000000000000000000000",
    726 => "10111110000100110110000000010111",
    727 => "00111111000011001010101111011000",
    728 => "00000000000000000000000000000000",
    729 => "00111111010101001001010001110100",
    730 => "00111110101111100111000001110010",
    731 => "10111110011010100111110011111001",
    732 => "00111111010001101101100000101000",
    733 => "00000000000000000000000000000000",
    734 => "00111111000111100101010111010110",
    735 => "00111111010000011110010111001101",
    736 => "00000000000000000000000000000000",
    737 => "10111110000100110110000000010000",
    738 => "00111111000011001010101111010101",
    739 => "00000000000000000000000000000000",
    740 => "00111111010101001001010001110110",
    741 => "00111110101111100111000001101111",
    742 => "10111110011010100111110011111100",
    743 => "00111111010001101101100000101000",
    744 => "00000000000000000000000000000000",
    745 => "00111111000111100101010111010110",
    746 => "00111111010000011110010111001011",
    747 => "00000000000000000000000000000000",
    748 => "10111110000100110110000000010000",
    749 => "00111111000011001010101111010101",
    750 => "00000000000000000000000000000000",
    751 => "00111111010101001001010001110110",
    752 => "00111111010000011110010111001011",
    753 => "00111111100100001000111100000001",
    754 => "00000000000000000000000000000000",
    755 => "00000000000000000000000000000000",
    756 => "00000000000000000000000000000000",
    757 => "00000000000000000000000000000000",
    758 => "10111111000000100111001000100111",
    759 => "10111110110000111110010100101100",
    760 => "00000000000000000000000000000000",
    761 => "00111111011011000100001010110101",
    762 => "00111100100011001000110111100000",
    763 => "00000000000000000000000000000000",
    764 => "10111110111111111110001011001010",
    765 => "00111111010000000101111101010111",
    766 => "00000000000000000000000000000000",
    767 => "00111111001001011000100111010100",
    768 => "00111110001001011010110100100111",
    769 => "10111110101100000110110001010100",
    770 => "10111110101010011010000001010011",
    771 => "00000000000000000000000000000000",
    772 => "00111111011100010110011010100000",
    773 => "00111101000001000011110110101010",
    774 => "00000000000000000000000000000000",
    775 => "10111110111101111101011010001000",
    776 => "00111111001111000111010011100010",
    777 => "00000000000000000000000000000000",
    778 => "00111111001010011001101110101000",
    779 => "00111110001010111001100011011001",
    780 => "10111110101011100000000100011001",
    781 => "10111110101010010010011101110101",
    782 => "00000000000000000000000000000000",
    783 => "00111111011100010111110000111100",
    784 => "00111101000001100101000101010111",
    785 => "00000000000000000000000000000000",
    786 => "10111110111101111000101000101000",
    787 => "00111111001111000101110001100011",
    788 => "00000000000000000000000000000000",
    789 => "00111111001010011011010001111000",
    790 => "00111110001010111110010111101110",
    791 => "10111110101011011110001000001001",
    792 => "10111110101010010010000101001000",
    793 => "00000000000000000000000000000000",
    794 => "00111111011100010111110101010111",
    795 => "00111101000001100110110000010111",
    796 => "00000000000000000000000000000000",
    797 => "10111110111101111000011001001111",
    798 => "00111111001111000101101100101100",
    799 => "00000000000000000000000000000000",
    800 => "00111111001010011011010110110010",
    801 => "00111110001010111110100111100000",
    802 => "10111110101011011110000001110001",
    803 => "10111110101010010010000011110111",
    804 => "00000000000000000000000000000000",
    805 => "00111111011100010111110101100101",
    806 => "00111101000001100110110101110110",
    807 => "00000000000000000000000000000000",
    808 => "10111110111101111000011000011011",
    809 => "00111111001111000101101100011011",
    810 => "00000000000000000000000000000000",
    811 => "00111111001010011011010111000011",
    812 => "00111101000001100110110101110110",
    813 => "00111110010011011000010101110000",
    814 => "00000000000000000000000000000000",
    815 => "00000000000000000000000000000000",
    816 => "00111111000110011001100110011010",
    817 => "00000000000000000000000000000000",
    818 => "00000000000000000000000000000000",
    819 => "10111111000000100111001000100111",
    820 => "00111111010010010010101101110110",
    821 => "00000000000000000000000000000000",
    822 => "00111111000110111001011010010100",
    823 => "00111110001011011110101101111011",
    824 => "00000000000000000000000000000000",
    825 => "10111110101011010001001010010101",
    826 => "00111111001101000100101010000010",
    827 => "00000000000000000000000000000000",
    828 => "00111111001100010010100000011001",
    829 => "00111110100010011101100100101001",
    830 => "10111110100011000001110111010000",
    831 => "00111111001011001100111111011110",
    832 => "00000000000000000000000000000000",
    833 => "00111111001110010011101011101110",
    834 => "00111110100111111110001101011101",
    835 => "00000000000000000000000000000000",
    836 => "10111110100000010111110011011100",
    837 => "00111111001010010111101100111010",
    838 => "00000000000000000000000000000000",
    839 => "00111111001111001001010011011100",
    840 => "00111110101001100010111100110110",
    841 => "10111110011111011000000001010110",
    842 => "00111111001010001000100101011101",
    843 => "00000000000000000000000000000000",
    844 => "00111111001111011000000110111110",
    845 => "00111110101001111011101001011111",
    846 => "00000000000000000000000000000000",
    847 => "10111110011111000011001000011110",
    848 => "00111111001010000100111001000011",
    849 => "00000000000000000000000000000000",
    850 => "00111111001111011011101100110100",
    851 => "00111110101010000001011101100000",
    852 => "10111110011110111110001111111101",
    853 => "00111111001010000100000001011100",
    854 => "00000000000000000000000000000000",
    855 => "00111111001111011100100010110010",
    856 => "00111110101010000010110100010000",
    857 => "00000000000000000000000000000000",
    858 => "10111110011110111101000111000101",
    859 => "00111111001010000011110100011111",
    860 => "00000000000000000000000000000000",
    861 => "00111111001111011100101111010110",
    862 => "00111110101010000011001000011010",
    863 => "10111110011110111100110110001100",
    864 => "00111111001010000011110001011100",
    865 => "00000000000000000000000000000000",
    866 => "00111111001111011100110010010010",
    867 => "00111110101010000011001101000010",
    868 => "00000000000000000000000000000000",
    869 => "10111110011110111100110010010011",
    870 => "00111111001010000011110000110010",
    871 => "00000000000000000000000000000000",
    872 => "00111111001111011100110010111100",
    873 => "00111110101010000011001101000010",
    874 => "00111111001010000011001101100110",
    875 => "00000000000000000000000000000000",
    876 => "00000000000000000000000000000000",
    877 => "00000000000000000000000000000000",
    878 => "00000000000000000000000000000000",
    879 => "00000000000000000000000000000000",
    880 => "00000000000000000000000000000000",
    881 => "00000000000000000000000000000000",
    882 => "10111111000000100111001000100111",
    883 => "10111111000110111001011100001010",
    884 => "00000000000000000000000000000000",
    885 => "00111111010010010010101100010100",
    886 => "00111101011100010010110000001100",
    887 => "00000000000000000000000000000000",
    888 => "10111110111001110101001110001000",
    889 => "00111111001110010000100001000000",
    890 => "00000000000000000000000000000000",
    891 => "00111111001011010000000100011111",
    892 => "00111110001111111001000001100110",
    893 => "10111110101001100100110001010000",
    894 => "10111111000001101110110000100000",
    895 => "00000000000000000000000000000000",
    896 => "00111111010110000111101110110101",
    897 => "00111101111000101010001111101111",
    898 => "00000000000000000000000000000000",
    899 => "10111110110010001101010000111000",
    900 => "00111111001101010101000110100101",
    901 => "00000000000000000000000000000000",
    902 => "00111111001100001000011100000000",
    903 => "00111110011010110010100001101100",
    904 => "10111110100101111001101111100010",
    905 => "10111111000001000010110100001101",
    906 => "00000000000000000000000000000000",
    907 => "00111111010110100100001010001010",
    908 => "00111101111101011110010010001110",
    909 => "00000000000000000000000000000000",
    910 => "10111110110000111110100011010010",
    911 => "00111111001101001010101101110111",
    912 => "00000000000000000000000000000000",
    913 => "00111111001100010010000001111100",
    914 => "00111110011100100110101001011000",
    915 => "10111110100101010110100110011100",
    916 => "10111111000000111011011000011001",
    917 => "00000000000000000000000000000000",
    918 => "00111111010110101000111000011010",
    919 => "00111101111110001100010111000001",
    920 => "00000000000000000000000000000000",
    921 => "10111110110000110011000011100010",
    922 => "00111111001101001001001001000000",
    923 => "00000000000000000000000000000000",
    924 => "00111111001100010011011110101011",
    925 => "00111110011100110111100110101111",
    926 => "10111110100101010001100011011100",
    927 => "10111111000000111010010010110011",
    928 => "00000000000000000000000000000000",
    929 => "00111111010110101001100100011110",
    930 => "00111101111110010010111110011100",
    931 => "00000000000000000000000000000000",
    932 => "10111110110000110001011010010010",
    933 => "00111111001101001000111010011110",
    934 => "00000000000000000000000000000000",
    935 => "00111111001100010011101100000001",
    936 => "00111101111110010010111110011100",
    937 => "00111110101110000001110000100001",
    938 => "00000000000000000000000000000000",
    939 => "00000000000000000000000000000000",
    940 => "00111110110011001100110011001110",
    941 => "00000000000000000000000000000000",
    942 => "00000000000000000000000000000000",
    943 => "10111111000000100111001000100111",
    944 => "00111111000110111001011100001100",
    945 => "00000000000000000000000000000000",
    946 => "00111111010010010010101100010010",
    947 => "00111101011100010010110000011000",
    948 => "00000000000000000000000000000000",
    949 => "10111110111001110101001110001000",
    950 => "00111111001110010000100001000000",
    951 => "00000000000000000000000000000000",
    952 => "00111111001011010000000100011111",
    953 => "00111110001111111001000001101000",
    954 => "10111110101001100100110001001111",
    955 => "00111111000001101110110000100010",
    956 => "00000000000000000000000000000000",
    957 => "00111111010110000111101110110100",
    958 => "00111101111000101010010000000001",
    959 => "00000000000000000000000000000000",
    960 => "10111110110010001101010000110101",
    961 => "00111111001101010101000110100011",
    962 => "00000000000000000000000000000000",
    963 => "00111111001100001000011100000010",
    964 => "00111110011010110010100001101010",
    965 => "10111110100101111001101111100101",
    966 => "00111111000001000010110100001111",
    967 => "00000000000000000000000000000000",
    968 => "00111111010110100100001010001001",
    969 => "00111101111101011110010010010001",
    970 => "00000000000000000000000000000000",
    971 => "10111110110000111110100011010010",
    972 => "00111111001101001010101101110111",
    973 => "00000000000000000000000000000000",
    974 => "00111111001100010010000001111100",
    975 => "00111110011100100110101001011000",
    976 => "10111110100101010110100110011100",
    977 => "00111111000000111011011000011010",
    978 => "00000000000000000000000000000000",
    979 => "00111111010110101000111000011001",
    980 => "00111101111110001100010111000001",
    981 => "00000000000000000000000000000000",
    982 => "10111110110000110011000011100010",
    983 => "00111111001101001001001001000000",
    984 => "00000000000000000000000000000000",
    985 => "00111111001100010011011110101011",
    986 => "00111110011100110111100110101111",
    987 => "10111110100101010001100011011100",
    988 => "00111111000000111010010010110101",
    989 => "00000000000000000000000000000000",
    990 => "00111111010110101001100100011101",
    991 => "00111101111110010010111110100100",
    992 => "00000000000000000000000000000000",
    993 => "10111110110000110001011010001111",
    994 => "00111111001101001000111010011110",
    995 => "00000000000000000000000000000000",
    996 => "00111111001100010011101100000001",
    997 => "00111101111110010010111110100100",
    998 => "00111110101110000001110000100110",
    999 => "00000000000000000000000000000000");

  constant b_lut : lut := (
    0 => "01000011000000000000000000000000",
    1 => "00000000000000000000000000000000",
    2 => "00111010001000100010010011101001",
    3 => "00111110101100101011011111111111",
    4 => "00111000001101010001111000111011",
    5 => "00111011010011010011011010110111",
    6 => "00111111000001100000100111111111",
    7 => "00111001101010111110101110110100",
    8 => "00111100001000100010101100010100",
    9 => "00111111010111110110010111111110",
    10 => "00111010101101010010011011011001",
    11 => "00111111010111110110010111111110",
    12 => "00111100001000100010101100010100",
    13 => "00111111010111110110010111111110",
    14 => "00111010101101010010011011011001",
    15 => "00000000000000000000000000000000",
    16 => "01000000000100000000000000000000",
    17 => "00111111100000000000000000000001",
    18 => "00000000000000000000000000000000",
    19 => "00111111100000000000000000000001",
    20 => "00000000000000000000000000000000",
    21 => "10111101110011001100110011001101",
    22 => "00000000000000000000000000000000",
    23 => "00111101110011001100110011001101",
    24 => "00111111011011011010000100000001",
    25 => "10110100101010111111000010010110",
    26 => "10111110000001100000101011000010",
    27 => "00110111010011010011101101011111",
    28 => "00111101110011001100110011001101",
    29 => "00111101110100000101100110000111",
    30 => "00111111011011011010000100000001",
    31 => "00111010100011101001010110000001",
    32 => "00111111100101011001101111100110",
    33 => "00111000101101110110100111011001",
    34 => "00111101110011001100110011001101",
    35 => "00111111011011011010000100000001",
    36 => "10110011010111010010110011111110",
    37 => "10111101101110100000000101011000",
    38 => "00110110001111100011111110101111",
    39 => "00111101110011001100110011001101",
    40 => "00111101110110000000111110000011",
    41 => "00111111011011011010000100000001",
    42 => "00111010101010010100000111001100",
    43 => "00111111100100110101101011101010",
    44 => "00111000111000110100001011111001",
    45 => "00111101110011001100110011001101",
    46 => "00111111011011011010000100000001",
    47 => "10110011011011111010011001001100",
    48 => "10111101101111010000001101111011",
    49 => "00110110010010101101101111000110",
    50 => "00111101110011001100110011001101",
    51 => "00111101110101111101101100100101",
    52 => "00111111011011011010000100000001",
    53 => "00111010101010001001001000000111",
    54 => "00111111100100110110100011100001",
    55 => "00111000111000100001110000011100",
    56 => "00111101110011001100110011001101",
    57 => "00111111011011011010000100000001",
    58 => "10110011011011110011100111000011",
    59 => "10111101101111001111001001011001",
    60 => "00110110010010101001001001000101",
    61 => "00111101110011001100110011001101",
    62 => "00111101110101111101110001010101",
    63 => "00111111011011011010000100000001",
    64 => "00111010101010001001010111100111",
    65 => "00111111100100110110100010010010",
    66 => "00111000111000100010001010011100",
    67 => "00111101110011001100110011001101",
    68 => "00111111011011011010000100000001",
    69 => "10110011011011110011110000110000",
    70 => "10111101101111001111001010111011",
    71 => "00110110010010101001001111101000",
    72 => "00111101110011001100110011001101",
    73 => "00111101110101111101110001001110",
    74 => "00111111011011011010000100000001",
    75 => "00111010101010001001010111011010",
    76 => "00111111100100110110100010010011",
    77 => "00111000111000100010001010000111",
    78 => "00111111000001111110100001010111",
    79 => "00111111100000000000000000000000",
    80 => "00111111110001001010010100100100",
    81 => "00111111100111101010011100000000",
    82 => "00000000000000000000000000000000",
    83 => "00111101110011001100110011001101",
    84 => "00111111011011011010000100000001",
    85 => "00111010100000011101110010001101",
    86 => "00111111100101101100110000011010",
    87 => "00111000101000110011000010011111",
    88 => "00111101110011001100110011001101",
    89 => "00111111001011101101000001000010",
    90 => "00111111011011011010000100000001",
    91 => "00111100011001010010111000000110",
    92 => "00111111010011110100000110101101",
    93 => "00111011000010111001000010001111",
    94 => "00111101110011001100110011001101",
    95 => "00111111011011011010000100000001",
    96 => "00111011000000011111100111011001",
    97 => "00111111010000000001110011100001",
    98 => "00111100010110000111111010000110",
    99 => "00111101110011001100110011001101",
    100 => "00111111010101110100101100101100",
    101 => "00111111011011011010000100000001",
    102 => "00111011000001010001110001101101",
    103 => "00111111010000010000011111100000",
    104 => "00111100010111001010100101101010",
    105 => "00111101110011001100110011001101",
    106 => "00111111011011011010000100000001",
    107 => "00111011000001001110010111001100",
    108 => "00111111010000001111100000000101",
    109 => "00111100010111000110000011110100",
    110 => "00111101110011001100110011001101",
    111 => "00111111010101110111100110010010",
    112 => "00111111011011011010000100000001",
    113 => "00111011000001001110100101101110",
    114 => "00111111010000001111100100010011",
    115 => "00111100010111000110010111000110",
    116 => "00111101110011001100110011001101",
    117 => "00111111011011011010000100000001",
    118 => "00111011000001001110100100101100",
    119 => "00111111010000001111100100000000",
    120 => "00111100010111000110010101101110",
    121 => "00111101110011001100110011001101",
    122 => "00111111010101110111100111000110",
    123 => "00111111011011011010000100000001",
    124 => "00111011000001001110100100110110",
    125 => "00111111010000001111100100000011",
    126 => "00111100010111000110010101111100",
    127 => "00111101110011001100110011001101",
    128 => "00111111011011011010000100000001",
    129 => "00111011000001001110100100101100",
    130 => "00111111010000001111100100000000",
    131 => "00111100010111000110010101101110",
    132 => "00111101110011001100110011001101",
    133 => "00111111010101110111100111000110",
    134 => "00111111011011011010000100000001",
    135 => "00111011000001001110100100110110",
    136 => "00111111010000001111100100000011",
    137 => "00111100010111000110010101111100",
    138 => "00111111001111011110000000110011",
    139 => "00111111100000000000000000000000",
    140 => "01000000000111101111000000011000",
    141 => "00111111110010011011011010000000",
    142 => "00000000000000000000000000000000",
    143 => "00111111011001100110011001101000",
    144 => "10111110100110011001100110011000",
    145 => "00000000000000000000000000000000",
    146 => "00111101110011001100110011001101",
    147 => "00111111011011011010000100000001",
    148 => "10111000101000110011010101011010",
    149 => "10111110110010010001000000100010",
    150 => "00111010100000011101111110010000",
    151 => "00111101110011001100110011001101",
    152 => "00111101111011111111000001000101",
    153 => "00111111011011011010000100000001",
    154 => "00111010111011111010001101000011",
    155 => "00111111100011100111101001000101",
    156 => "00111001001011110111110111100011",
    157 => "00111101110011001100110011001101",
    158 => "00111111011011011010000100000001",
    159 => "10110111100000000010111110010101",
    160 => "10111110100100010011000011100110",
    161 => "00111001100011010100000111001011",
    162 => "00111101110011001100110011001101",
    163 => "00111110000110010001011110000011",
    164 => "00111111011011011010000100000001",
    165 => "00111011001011011011111011010111",
    166 => "00111111100010001100011000101111",
    167 => "00111001100010111001111111101010",
    168 => "00111101110011001100110011001101",
    169 => "00111111011011011010000100000001",
    170 => "10110111011110000010001110011100",
    171 => "10111110100100000011111100001111",
    172 => "00111001100010011001110111001001",
    173 => "00111101110011001100110011001101",
    174 => "00111110000110010111111000010110",
    175 => "00111111011011011010000100000001",
    176 => "00111011001011100010011010011010",
    177 => "00111111100010001011110010011000",
    178 => "00111001100011000000100000101100",
    179 => "00111101110011001100110011001101",
    180 => "00111111011011011010000100000001",
    181 => "10110111011101111100000100101011",
    182 => "10111110100100000011001110011011",
    183 => "00111001100010010111001000011001",
    184 => "00111101110011001100110011001101",
    185 => "00111110000110011000001011100110",
    186 => "00111111011011011010000100000001",
    187 => "00111011001011100010101101111001",
    188 => "00111111100010001011110000100101",
    189 => "00111001100011000000110100001111",
    190 => "00111101110011001100110011001101",
    191 => "00111111011011011010000100000001",
    192 => "10110111011101111011110010011100",
    193 => "10111110100100000011001100010011",
    194 => "00111001100010010111000000010011",
    195 => "00111101110011001100110011001101",
    196 => "00111110000110011000001100100000",
    197 => "00111111011011011010000100000001",
    198 => "00111011001011100010101110101110",
    199 => "00111111100010001011110000100000",
    200 => "00111001100011000000110101000110",
    201 => "00111110111111100001011000010011",
    202 => "00111111100000000000000000000000",
    203 => "00111111110001011110100100011100",
    204 => "00111111100111110010100101111011",
    205 => "00111101110011001100110011001101",
    206 => "00000000000000000000000000000000",
    207 => "00111101110011001100110011001101",
    208 => "00111111011011011010000100000001",
    209 => "00111011111110101000001101110001",
    210 => "00111111011010101001001011010101",
    211 => "00111010100000110010101110101011",
    212 => "00111101110011001100110011001101",
    213 => "00111110100010100010100011110001",
    214 => "00111111011011011010000100000001",
    215 => "00111011100001111110110100101110",
    216 => "00111111100000010010100101000010",
    217 => "00111001111101000101011000010011",
    218 => "00111101110011001100110011001101",
    219 => "00111111011011011010000100000001",
    220 => "00111010001011000111011110101000",
    221 => "00111111000110100001000101111000",
    222 => "00111011101100110001101001110000",
    223 => "00111101110011001100110011001101",
    224 => "00111110111011111110010110110110",
    225 => "00111111011011011010000100000001",
    226 => "00111100000001101011101100101001",
    227 => "00111111011001110111110111000110",
    228 => "00111010100011111011000000010101",
    229 => "00111101110011001100110011001101",
    230 => "00111111011011011010000100000001",
    231 => "00111010000100100111011000100100",
    232 => "00111111000101010001110100000001",
    233 => "00111011100111010010011010011001",
    234 => "00111101110011001100110011001101",
    235 => "00111110111100011010001010100000",
    236 => "00111111011011011010000100000001",
    237 => "00111100000010000001101001111110",
    238 => "00111111011001110000111011110101",
    239 => "00111010100100011000010100001011",
    240 => "00111101110011001100110011001101",
    241 => "00111111011011011010000100000001",
    242 => "00111010000100100110011010001010",
    243 => "00111111000101010001100111010100",
    244 => "00111011100111010001100100110111",
    245 => "00111101110011001100110011001101",
    246 => "00111110111100011010001110011000",
    247 => "00111111011011011010000100000001",
    248 => "00111100000010000001101100111010",
    249 => "00111111011001110000111010111010",
    250 => "00111010100100011000011000000110",
    251 => "00111101110011001100110011001101",
    252 => "00111111011011011010000100000001",
    253 => "00111010000100100110011001111011",
    254 => "00111111000101010001100111010001",
    255 => "00111011100111010001100100101010",
    256 => "00111101110011001100110011001101",
    257 => "00111110111100011010001110100101",
    258 => "00111111011011011010000100000001",
    259 => "00111100000010000001101101000111",
    260 => "00111111011001110000111010110110",
    261 => "00111010100100011000011000011000",
    262 => "00111111010000011110010111001101",
    263 => "00111111100000000000000000000000",
    264 => "01000000000010000100011110000010",
    265 => "00111111101110101100100000101111",
    266 => "00000000000000000000000000000000",
    267 => "00111101110011001100110011001101",
    268 => "00111111011011011010000100000001",
    269 => "10111010100000110010110111110111",
    270 => "10111111001001111000110101110001",
    271 => "00111011111110101000011011101111",
    272 => "00111101110011001100110011001101",
    273 => "00111110001000101011000101101010",
    274 => "00111111011011011010000100000001",
    275 => "00111011001101101010000110010101",
    276 => "00111111100001111111011110101111",
    277 => "00111001100101001001101101011011",
    278 => "00111101110011001100110011001101",
    279 => "00111111011011011010000100000001",
    280 => "10111001001111111011001001111001",
    281 => "10111110111011101000001101110000",
    282 => "00111011000000001001011101101110",
    283 => "00111101110011001100110011001101",
    284 => "00111110100000100100111001000101",
    285 => "00111111011011011010000100000001",
    286 => "00111011100000001001010110111001",
    287 => "00111111100000100010011100000000",
    288 => "00111001111000111111001111101101",
    289 => "00111101110011001100110011001101",
    290 => "00111111011011011010000100000001",
    291 => "10111001000001001111101011010010",
    292 => "10111110110111011011000010111100",
    293 => "00111010101111111111001000011000",
    294 => "00111101110011001100110011001101",
    295 => "00111110100001101110011001010010",
    296 => "00111111011011011010000100000001",
    297 => "00111011100001001101000011011110",
    298 => "00111111100000011001001101111011",
    299 => "00111001111011010101110111101111",
    300 => "00111101110011001100110011001101",
    301 => "00111111011011011010000100000001",
    302 => "10111001000000100001110011101011",
    303 => "10111110110111001011100111100110",
    304 => "00111010101111001010000011001001",
    305 => "00111101110011001100110011001101",
    306 => "00111110100001110010000111000011",
    307 => "00111111011011011010000100000001",
    308 => "00111011100001010000100011010000",
    309 => "00111111100000011000101111110101",
    310 => "00111001111011011101101011110001",
    311 => "00111101110011001100110011001101",
    312 => "00111111011011011010000100000001",
    313 => "10111001000000011111100111101111",
    314 => "10111110110111001010111000000110",
    315 => "00111010101111000111100000110100",
    316 => "00111101110011001100110011001101",
    317 => "00111110100001110010010010010110",
    318 => "00111111011011011010000100000001",
    319 => "00111011100001010000101101110101",
    320 => "00111111100000011000101110011010",
    321 => "00111001111011011110000011011101",
    322 => "00111111001011001110001101000010",
    323 => "00111111100000000000000000000000",
    324 => "00111111111010110110110111111010",
    325 => "00111111101011011001100000100101",
    326 => "00111101110011001100110011001101",
    327 => "00000000000000000000000000000000",
    328 => "00111101110011001100110011001101",
    329 => "00111111011011011010000100000001",
    330 => "00111010100000110010111000000010",
    331 => "00111111001001111000110101110100",
    332 => "00111011111110101000011100000100",
    333 => "00111101110011001100110011001101",
    334 => "00111110001000101011000101101100",
    335 => "00111111011011011010000100000001",
    336 => "00111011001101101010000110010101",
    337 => "00111111100001111111011110101111",
    338 => "00111001100101001001101101011011",
    339 => "00111101110011001100110011001101",
    340 => "00111111011011011010000100000001",
    341 => "00111001001111111011001010000101",
    342 => "00111110111011101000001101110011",
    343 => "00111011000000001001011101110101",
    344 => "00111101110011001100110011001101",
    345 => "00111110100000100100111001001001",
    346 => "00111111011011011010000100000001",
    347 => "00111011100000001001010111000001",
    348 => "00111111100000100010011011111111",
    349 => "00111001111000111111001111111110",
    350 => "00111101110011001100110011001101",
    351 => "00111111011011011010000100000001",
    352 => "00111001000001001111101011011100",
    353 => "00111110110111011011000010111111",
    354 => "00111010101111111111001000100011",
    355 => "00111101110011001100110011001101",
    356 => "00111110100001101110011001010011",
    357 => "00111111011011011010000100000001",
    358 => "00111011100001001101000011010110",
    359 => "00111111100000011001001101111100",
    360 => "00111001111011010101110111011111",
    361 => "00111101110011001100110011001101",
    362 => "00111111011011011010000100000001",
    363 => "00111001000000100001110011101111",
    364 => "00111110110111001011100111100111",
    365 => "00111010101111001010000011001101",
    366 => "00111101110011001100110011001101",
    367 => "00111110100001110010000111001001",
    368 => "00111111011011011010000100000001",
    369 => "00111011100001010000100011011000",
    370 => "00111111100000011000101111110100",
    371 => "00111001111011011101101100000001",
    372 => "00111101110011001100110011001101",
    373 => "00111111011011011010000100000001",
    374 => "00111001000000011111100111111001",
    375 => "00111110110111001010111000001001",
    376 => "00111010101111000111100000111110",
    377 => "00111101110011001100110011001101",
    378 => "00111110100001110010010010011001",
    379 => "00111111011011011010000100000001",
    380 => "00111011100001010000101101110101",
    381 => "00111111100000011000101110011010",
    382 => "00111001111011011110000011011101",
    383 => "00111111001011001110001101000111",
    384 => "00111111100000000000000000000000",
    385 => "00111111111010110110110111111101",
    386 => "00111111101011011001100000100110",
    387 => "00000000000000000000000000000000",
    388 => "00111111011001100110011001101000",
    389 => "10111111001100110011001100110010",
    390 => "00000000000000000000000000000000",
    391 => "00111101110011001100110011001101",
    392 => "00111111011011011010000100000001",
    393 => "10111011101100000110000011111101",
    394 => "10111111011010101001001011010011",
    395 => "00111100111100001001101100111010",
    396 => "00111101110011001100110011001101",
    397 => "00111110100010100010100100010100",
    398 => "00111111011011011010000100000001",
    399 => "00111011100001111110110101001110",
    400 => "00111111100000010010100100111110",
    401 => "00111001111101000101011001011001",
    402 => "00111101110011001100110011001101",
    403 => "00111111011011011010000100000001",
    404 => "10111010001011000111011110001000",
    405 => "10111111000110100001000101110010",
    406 => "00111011101100110001101001010100",
    407 => "00111101110011001100110011001101",
    408 => "00111110111011111110010110111101",
    409 => "00111111011011011010000100000001",
    410 => "00111100000001101011101100101110",
    411 => "00111111011001110111110111000100",
    412 => "00111010100011111011000000011101",
    413 => "00111101110011001100110011001101",
    414 => "00111111011011011010000100000001",
    415 => "10111010000100100111011000011001",
    416 => "10111111000101010001110011111111",
    417 => "00111011100111010010011010010001",
    418 => "00111101110011001100110011001101",
    419 => "00111110111100011010001010010110",
    420 => "00111111011011011010000100000001",
    421 => "00111100000010000001101001110010",
    422 => "00111111011001110000111011111001",
    423 => "00111010100100011000010011111010",
    424 => "00111101110011001100110011001101",
    425 => "00111111011011011010000100000001",
    426 => "10111010000100100110011010000000",
    427 => "10111111000101010001100111010010",
    428 => "00111011100111010001100100101110",
    429 => "00111101110011001100110011001101",
    430 => "00111110111100011010001110011101",
    431 => "00111111011011011010000100000001",
    432 => "00111100000010000001101101000111",
    433 => "00111111011001110000111010110110",
    434 => "00111010100100011000011000011000",
    435 => "00111101110011001100110011001101",
    436 => "00111111011011011010000100000001",
    437 => "10111010000100100110011010000000",
    438 => "10111111000101010001100111010010",
    439 => "00111011100111010001100100101110",
    440 => "00111101110011001100110011001101",
    441 => "00111110111100011010001110011101",
    442 => "00111111011011011010000100000001",
    443 => "00111100000010000001101101000111",
    444 => "00111111011001110000111010110110",
    445 => "00111010100100011000011000011000",
    446 => "00111111010000011110010111001000",
    447 => "00111111100000000000000000000000",
    448 => "01000000000010000100011101111111",
    449 => "00111111101110101100100000101101",
    450 => "00111101110011001100110011001101",
    451 => "00000000000000000000000000000000",
    452 => "00111101110011001100110011001101",
    453 => "00111111011011011010000100000001",
    454 => "00111000101000110011010101100000",
    455 => "00111110110010010001000000100100",
    456 => "00111010100000011101111110010101",
    457 => "00111101110011001100110011001101",
    458 => "00111101111011111111000001000110",
    459 => "00111111011011011010000100000001",
    460 => "00111010111011111010001101000011",
    461 => "00111111100011100111101001000101",
    462 => "00111001001011110111110111100011",
    463 => "00111101110011001100110011001101",
    464 => "00111111011011011010000100000001",
    465 => "00110111100000000010111110011110",
    466 => "00111110100100010011000011101000",
    467 => "00111001100011010100000111010010",
    468 => "00111101110011001100110011001101",
    469 => "00111110000110010001011110000100",
    470 => "00111111011011011010000100000001",
    471 => "00111011001011011011111011010111",
    472 => "00111111100010001100011000101111",
    473 => "00111001100010111001111111101010",
    474 => "00111101110011001100110011001101",
    475 => "00111111011011011010000100000001",
    476 => "00110111011110000010001110101111",
    477 => "00111110100100000011111100010001",
    478 => "00111001100010011001110111010000",
    479 => "00111101110011001100110011001101",
    480 => "00111110000110010111111000011000",
    481 => "00111111011011011010000100000001",
    482 => "00111011001011100010011010011010",
    483 => "00111111100010001011110010011000",
    484 => "00111001100011000000100000101100",
    485 => "00111101110011001100110011001101",
    486 => "00111111011011011010000100000001",
    487 => "00110111011101111100000100111110",
    488 => "00111110100100000011001110011101",
    489 => "00111001100010010111001000100001",
    490 => "00111101110011001100110011001101",
    491 => "00111110000110011000001011101000",
    492 => "00111111011011011010000100000001",
    493 => "00111011001011100010101101111001",
    494 => "00111111100010001011110000100101",
    495 => "00111001100011000000110100001111",
    496 => "00111101110011001100110011001101",
    497 => "00111111011011011010000100000001",
    498 => "00110111011101111011110010101100",
    499 => "00111110100100000011001100010101",
    500 => "00111001100010010111000000011011",
    501 => "00111101110011001100110011001101",
    502 => "00111110000110011000001100100010",
    503 => "00111111011011011010000100000001",
    504 => "00111011001011100010101110111001",
    505 => "00111111100010001011110000011111",
    506 => "00111001100011000000110101010010",
    507 => "00111110111111100001011000011001",
    508 => "00111111100000000000000000000000",
    509 => "00111111110001011110100100011110",
    510 => "00111111100111110010100101111011",
    511 => "00000000000000000000000000000000",
    512 => "00111101110011001100110011001101",
    513 => "00111111011011011010000100000001",
    514 => "10111100100110101110101110100110",
    515 => "10111111100101101100110000011010",
    516 => "00111101101001000101111011110101",
    517 => "00111101110011001100110011001101",
    518 => "00111111001011101101100011000110",
    519 => "00111111011011011010000100000001",
    520 => "00111100011001010011110101110110",
    521 => "00111111010011110011111001100101",
    522 => "00111011000010111001110001010001",
    523 => "00111101110011001100110011001101",
    524 => "00111111011011011010000100000001",
    525 => "10111011000000011111101001100101",
    526 => "10111111010000000001110100001010",
    527 => "00111100010110000111111100111111",
    528 => "00111101110011001100110011001101",
    529 => "00111111010101110100101100110000",
    530 => "00111111011011011010000100000001",
    531 => "00111011000001010001110001100111",
    532 => "00111111010000010000011111011110",
    533 => "00111100010111001010100101100000",
    534 => "00111101110011001100110011001101",
    535 => "00111111011011011010000100000001",
    536 => "10111011000001001110010111001100",
    537 => "10111111010000001111100000000101",
    538 => "00111100010111000110000011110100",
    539 => "00111101110011001100110011001101",
    540 => "00111111010101110111100110001110",
    541 => "00111111011011011010000100000001",
    542 => "00111011000001001110100101110101",
    543 => "00111111010000001111100100010101",
    544 => "00111100010111000110010111001110",
    545 => "00111101110011001100110011001101",
    546 => "00111111011011011010000100000001",
    547 => "10111011000001001110100100010111",
    548 => "10111111010000001111100011111010",
    549 => "00111100010111000110010101010100",
    550 => "00111101110011001100110011001101",
    551 => "00111111010101110111100110111100",
    552 => "00111111011011011010000100000001",
    553 => "00111011000001001110100100111101",
    554 => "00111111010000001111100100000101",
    555 => "00111100010111000110010110000110",
    556 => "00111101110011001100110011001101",
    557 => "00111111011011011010000100000001",
    558 => "10111011000001001110100100110000",
    559 => "10111111010000001111100100000001",
    560 => "00111100010111000110010101110100",
    561 => "00111101110011001100110011001101",
    562 => "00111111010101110111100111000100",
    563 => "00111111011011011010000100000001",
    564 => "00111011000001001110100100110110",
    565 => "00111111010000001111100100000011",
    566 => "00111100010111000110010101111100",
    567 => "00111111001111011110000000110001",
    568 => "00111111100000000000000000000000",
    569 => "01000000000111101111000000010111",
    570 => "00111111110010011011011001111111",
    571 => "00111101110011001100110011001101",
    572 => "00000000000000000000000000000000",
    573 => "00111101110011001100110011001101",
    574 => "00111111011011011010000100000001",
    575 => "00110100101010111111000010010110",
    576 => "00111110000001100000101011000010",
    577 => "00110111010011010011101101011111",
    578 => "00111101110011001100110011001101",
    579 => "00111101110100000101100110000111",
    580 => "00111111011011011010000100000001",
    581 => "00111010100011101001010110000001",
    582 => "00111111100101011001101111100110",
    583 => "00111000101101110110100111011001",
    584 => "00111101110011001100110011001101",
    585 => "00111111011011011010000100000001",
    586 => "00110011010111010010110011111110",
    587 => "00111101101110100000000101011000",
    588 => "00110110001111100011111110101111",
    589 => "00111101110011001100110011001101",
    590 => "00111101110110000000111110000011",
    591 => "00111111011011011010000100000001",
    592 => "00111010101010010100000111001100",
    593 => "00111111100100110101101011101010",
    594 => "00111000111000110100001011111001",
    595 => "00111101110011001100110011001101",
    596 => "00111111011011011010000100000001",
    597 => "00110011011011111010011001001100",
    598 => "00111101101111010000001101111011",
    599 => "00110110010010101101101111000110",
    600 => "00111101110011001100110011001101",
    601 => "00111101110101111101101100100101",
    602 => "00111111011011011010000100000001",
    603 => "00111010101010001001001000000111",
    604 => "00111111100100110110100011100001",
    605 => "00111000111000100001110000011100",
    606 => "00111101110011001100110011001101",
    607 => "00111111011011011010000100000001",
    608 => "00110011011011110011100111000011",
    609 => "00111101101111001111001001011001",
    610 => "00110110010010101001001001000101",
    611 => "00111101110011001100110011001101",
    612 => "00111101110101111101110001010101",
    613 => "00111111011011011010000100000001",
    614 => "00111010101010001001010111100111",
    615 => "00111111100100110110100010010010",
    616 => "00111000111000100010001010011100",
    617 => "00111101110011001100110011001101",
    618 => "00111111011011011010000100000001",
    619 => "00110011011011110011110000110000",
    620 => "00111101101111001111001010111011",
    621 => "00110110010010101001001111101000",
    622 => "00111101110011001100110011001101",
    623 => "00111101110101111101110001001110",
    624 => "00111111011011011010000100000001",
    625 => "00111010101010001001010111011010",
    626 => "00111111100100110110100010010011",
    627 => "00111000111000100010001010000111",
    628 => "00111111000001111110100001010111",
    629 => "00111111100000000000000000000000",
    630 => "00111111110001001010010100100100",
    631 => "00111111100111101010011100000000",
    632 => "00000000000000000000000000000000",
    633 => "00111111001100110011001100110110",
    634 => "10111101110011001100110011000000",
    635 => "00000000000000000000000000000000",
    636 => "00111101110011001100110011001101",
    637 => "00111111011011011010000100000001",
    638 => "10110100101010111111000001100100",
    639 => "10111110000001100000101010111010",
    640 => "00110111010011010011101100101110",
    641 => "00111101110011001100110011001101",
    642 => "00111101110100000101100110000110",
    643 => "00111111011011011010000100000001",
    644 => "00111100000000101110000001010111",
    645 => "00111111011010001011100110100000",
    646 => "00111010100010101001000101001100",
    647 => "00111101110011001100110011001101",
    648 => "00111111011011011010000100000001",
    649 => "10110100000111110110001001001000",
    650 => "10111101111001011101111000111000",
    651 => "00110110110111011101111110011110",
    652 => "00111101110011001100110011001101",
    653 => "00111101110100111100001111110001",
    654 => "00111111011011011010000100000001",
    655 => "00111100000001111111111110101010",
    656 => "00111111011001110001011101100100",
    657 => "00111010100100010110000100110001",
    658 => "00111101110011001100110011001101",
    659 => "00111111011011011010000100000001",
    660 => "10110100001000000000111010101110",
    661 => "10111101111001100000111111011101",
    662 => "00110110110111101001111110000110",
    663 => "00111101110011001100110011001101",
    664 => "00111101110100111011101111010000",
    665 => "00111111011011011010000100000001",
    666 => "00111100000001111111001111001001",
    667 => "00111111011001110001101100100000",
    668 => "00111010100100010101000101010001",
    669 => "00111101110011001100110011001101",
    670 => "00111111011011011010000100000001",
    671 => "10110100001000000000110100111101",
    672 => "10111101111001100000111101110011",
    673 => "00110110110111101001110111101101",
    674 => "00111101110011001100110011001101",
    675 => "00111101110100111011101111100010",
    676 => "00111111011011011010000100000001",
    677 => "00111100000001111111001111100000",
    678 => "00111111011001110001101100011001",
    679 => "00111010100100010101000101101110",
    680 => "00111101110011001100110011001101",
    681 => "00111111011011011010000100000001",
    682 => "10110100001000000000110100111101",
    683 => "10111101111001100000111101110011",
    684 => "00110110110111101001110111101101",
    685 => "00111101110011001100110011001101",
    686 => "00111101110100111011101111100010",
    687 => "00111111011011011010000100000001",
    688 => "00111100000001111111001111100000",
    689 => "00111111011001110001101100011001",
    690 => "00111010100100010101000101101110",
    691 => "00111110001010100000100001110010",
    692 => "00111111100000000000000000000000",
    693 => "00111111100101011011000000000000",
    694 => "00111111100010100110101101101110",
    695 => "00111101110011001100110011001101",
    696 => "00000000000000000000000000000000",
    697 => "00111101110011001100110011001101",
    698 => "00111111011011011010000100000001",
    699 => "00111010100000011101110010000011",
    700 => "00111111100101101100110000011011",
    701 => "00111000101000110011000010001110",
    702 => "00111101110011001100110011001101",
    703 => "00111111001011101101000001001000",
    704 => "00111111011011011010000100000001",
    705 => "00111010010110000100000010001000",
    706 => "00111111001000010011001100010100",
    707 => "00111011110101101010001101000011",
    708 => "00111101110011001100110011001101",
    709 => "00111111011011011010000100000001",
    710 => "00111100000001000101000010011011",
    711 => "00111111011010000100001011110011",
    712 => "00111010100011000111100101011001",
    713 => "00111101110011001100110011001101",
    714 => "00111111010110110101100001111000",
    715 => "00111111011011011010000100000001",
    716 => "00111010000100101001010100011011",
    717 => "00111111000101010010001101001111",
    718 => "00111011100111010100000100101110",
    719 => "00111101110011001100110011001101",
    720 => "00111111011011011010000100000001",
    721 => "00111100000010000001100011010101",
    722 => "00111111011001110000111101111011",
    723 => "00111010100100011000001011010010",
    724 => "00111101110011001100110011001101",
    725 => "00111111010110110111111101010110",
    726 => "00111111011011011010000100000001",
    727 => "00111010000100100110011010011010",
    728 => "00111111000101010001100111010111",
    729 => "00111011100111010001100101000011",
    730 => "00111101110011001100110011001101",
    731 => "00111111011011011010000100000001",
    732 => "00111100000010000001101101000111",
    733 => "00111111011001110000111010110110",
    734 => "00111010100100011000011000011000",
    735 => "00111101110011001100110011001101",
    736 => "00111111010110110111111101100110",
    737 => "00111111011011011010000100000001",
    738 => "00111010000100100110011010001010",
    739 => "00111111000101010001100111010100",
    740 => "00111011100111010001100100110111",
    741 => "00111101110011001100110011001101",
    742 => "00111111011011011010000100000001",
    743 => "00111100000010000001101101000111",
    744 => "00111111011001110000111010110110",
    745 => "00111010100100011000011000011000",
    746 => "00111101110011001100110011001101",
    747 => "00111111010110110111111101100100",
    748 => "00111111011011011010000100000001",
    749 => "00111010000100100110011010001010",
    750 => "00111111000101010001100111010100",
    751 => "00111011100111010001100100110111",
    752 => "00111110101111100111000001101111",
    753 => "00111111100000000000000000000000",
    754 => "01000000000010000100011110000000",
    755 => "00111111101110101100100000101110",
    756 => "00000000000000000000000000000000",
    757 => "00111101110011001100110011001101",
    758 => "00111111011011011010000100000001",
    759 => "10111000101000110011010101011010",
    760 => "10111110110010010001000000100010",
    761 => "00111010100000011101111110010000",
    762 => "00111101110011001100110011001101",
    763 => "00111101111011111111000001000101",
    764 => "00111111011011011010000100000001",
    765 => "00111100001010001010110011100110",
    766 => "00111111010111011010000111000100",
    767 => "00111010101111100100100001101111",
    768 => "00111101110011001100110011001101",
    769 => "00111111011011011010000100000001",
    770 => "10111000000110011000110100001011",
    771 => "10111110101011001110100111001001",
    772 => "00111010000011100001010010001110",
    773 => "00111101110011001100110011001101",
    774 => "00111110000001110111010111010001",
    775 => "00111111011011011010000100000001",
    776 => "00111100001111100001001101101111",
    777 => "00111111010110000010100100101010",
    778 => "00111010110111001110110010110001",
    779 => "00111101110011001100110011001101",
    780 => "00111111011011011010000100000001",
    781 => "10111000000101110101011101010010",
    782 => "10111110101011000110100110100010",
    783 => "00111010000011000111000100101110",
    784 => "00111101110011001100110011001101",
    785 => "00111110000001111111101010111100",
    786 => "00111111011011011010000100000001",
    787 => "00111100001111101001110101100111",
    788 => "00111111010110000000011101110100",
    789 => "00111010110111011011010100111000",
    790 => "00111101110011001100110011001101",
    791 => "00111111011011011010000100000001",
    792 => "10111000000101110011101010010011",
    793 => "10111110101011000110001100010101",
    794 => "00111010000011000101101111010111",
    795 => "00111101110011001100110011001101",
    796 => "00111110000010000000000101101100",
    797 => "00111111011011011010000100000001",
    798 => "00111100001111101010010001000001",
    799 => "00111111010110000000010111001000",
    800 => "00111010110111011011111100101101",
    801 => "00111101110011001100110011001101",
    802 => "00111111011011011010000100000001",
    803 => "10111000000101110011100100011111",
    804 => "10111110101011000110001011000000",
    805 => "00111010000011000101101011000010",
    806 => "00111101110011001100110011001101",
    807 => "00111110000010000000000111000100",
    808 => "00111111011011011010000100000001",
    809 => "00111100001111101010010010011111",
    810 => "00111111010110000000010110110001",
    811 => "00111010110111011011111110110101",
    812 => "00111110001010111110101000010011",
    813 => "00111111100000000000000000000000",
    814 => "00111111100110011011000010101110",
    815 => "00111111100011000100001000010100",
    816 => "00111101110011001100110011001101",
    817 => "00000000000000000000000000000000",
    818 => "00111101110011001100110011001101",
    819 => "00111111011011011010000100000001",
    820 => "00111011111110101000001101110001",
    821 => "00111111011010101001001011010101",
    822 => "00111010100000110010101110101011",
    823 => "00111101110011001100110011001101",
    824 => "00111110100010100010100011110001",
    825 => "00111111011011011010000100000001",
    826 => "00111011001000101001111001000110",
    827 => "00111111010010001110101011011011",
    828 => "00111100100000010111111101011010",
    829 => "00111101110011001100110011001101",
    830 => "00111111011011011010000100000001",
    831 => "00111010111110000100001010000011",
    832 => "00111111001111100101101001001001",
    833 => "00111100010100001010101100100101",
    834 => "00111101110011001100110011001101",
    835 => "00111110110100110001011010010000",
    836 => "00111111011011011010000100000001",
    837 => "00111010110110111110011110010110",
    838 => "00111111001110011100101001111100",
    839 => "00111100001111010101111110100001",
    840 => "00111101110011001100110011001101",
    841 => "00111111011011011010000100000001",
    842 => "00111010110101000110111111001000",
    843 => "00111111001110001000001011110110",
    844 => "00111100001110000011011000000000",
    845 => "00111101110011001100110011001101",
    846 => "00111110110110101110110110010010",
    847 => "00111111011011011010000100000001",
    848 => "00111010110100101010010111111110",
    849 => "00111111001110000011001100101011",
    850 => "00111100001101101111100000100111",
    851 => "00111101110011001100110011001101",
    852 => "00111111011011011010000100000001",
    853 => "00111010110100100011101011010001",
    854 => "00111111001110000010000001101001",
    855 => "00111100001101101010110110101011",
    856 => "00111101110011001100110011001101",
    857 => "00111110110110110110000001000011",
    858 => "00111111011011011010000100000001",
    859 => "00111010110100100010000111100100",
    860 => "00111111001110000001110000001011",
    861 => "00111100001101101001110001010111",
    862 => "00111101110011001100110011001101",
    863 => "00111111011011011010000100000001",
    864 => "00111010110100100001110000001110",
    865 => "00111111001110000001101100000101",
    866 => "00111100001101101001100001001001",
    867 => "00111101110011001100110011001101",
    868 => "00111110110110110110011001110101",
    869 => "00111111011011011010000100000001",
    870 => "00111010110100100001101011000001",
    871 => "00111111001110000001101011001011",
    872 => "00111100001101101001011101100010",
    873 => "00111110101010000011001110001011",
    874 => "00111111100000000000000000000000",
    875 => "00111111110101000001100110110011",
    876 => "00111111101001001100010011100010",
    877 => "00000000000000000000000000000000",
    878 => "00111111001100110011001100110110",
    879 => "10111110111111111111111111111110",
    880 => "00000000000000000000000000000000",
    881 => "00111101110011001100110011001101",
    882 => "00111111011011011010000100000001",
    883 => "10111010100000110010110111110111",
    884 => "10111111001001111000110101110001",
    885 => "00111011111110101000011011101111",
    886 => "00111101110011001100110011001101",
    887 => "00111110001000101011000101101010",
    888 => "00111111011011011010000100000001",
    889 => "00111100010100011101011001101000",
    890 => "00111111010100111000000101001100",
    891 => "00111010111110011111111111011110",
    892 => "00111101110011001100110011001101",
    893 => "00111111011011011010000100000001",
    894 => "10111001111001110101110110111100",
    895 => "10111111000011100011110111000101",
    896 => "00111011100000100001111101110110",
    897 => "00111101110011001100110011001101",
    898 => "00111110010101111011100001011110",
    899 => "00111111011011011010000100000001",
    900 => "00111100011010000101111011111100",
    901 => "00111111010011101001010011101010",
    902 => "00111011000011011111111110000110",
    903 => "00111101110011001100110011001101",
    904 => "00111111011011011010000100000001",
    905 => "10111001110011100011101100001111",
    906 => "10111111000010110000000111000100",
    907 => "00111011011011010101111011001111",
    908 => "00111101110011001100110011001101",
    909 => "00111110011000010101100010101110",
    910 => "00111111011011011010000100000001",
    911 => "00111100011011000110110110100000",
    912 => "00111111010011011011101111010011",
    913 => "00111011000100010001101010100000",
    914 => "00111101110011001100110011001101",
    915 => "00111111011011011010000100000001",
    916 => "10111001110010100011100011010101",
    917 => "10111111000010100111011001010110",
    918 => "00111011011010011010110000000101",
    919 => "00111101110011001100110011001101",
    920 => "00111110011000101100100101000111",
    921 => "00111111011011011010000100000001",
    922 => "00111100011011010000110000000011",
    923 => "00111111010011011001101011110111",
    924 => "00111011000100011001010000101011",
    925 => "00111101110011001100110011001101",
    926 => "00111111011011011010000100000001",
    927 => "10111001110010011010010000111000",
    928 => "10111111000010100110000111110110",
    929 => "00111011011010010010001010011001",
    930 => "00111101110011001100110011001101",
    931 => "00111110011000101111111000110100",
    932 => "00111111011011011010000100000001",
    933 => "00111100011011010010001011011001",
    934 => "00111111010011011001011000111100",
    935 => "00111011000100011010010110110010",
    936 => "00111110011100111010000001110100",
    937 => "00111111100000000000000000000000",
    938 => "00111111101011100000011100001000",
    939 => "00111111100101010011111111110101",
    940 => "00111101110011001100110011001101",
    941 => "00000000000000000000000000000000",
    942 => "00111101110011001100110011001101",
    943 => "00111111011011011010000100000001",
    944 => "00111010100000110010111000000010",
    945 => "00111111001001111000110101110100",
    946 => "00111011111110101000011100000100",
    947 => "00111101110011001100110011001101",
    948 => "00111110001000101011000101101100",
    949 => "00111111011011011010000100000001",
    950 => "00111100010100011101011001101000",
    951 => "00111111010100111000000101001100",
    952 => "00111010111110011111111111011110",
    953 => "00111101110011001100110011001101",
    954 => "00111111011011011010000100000001",
    955 => "00111001111001110101110111001101",
    956 => "00111111000011100011110111000111",
    957 => "00111011100000100001111101111110",
    958 => "00111101110011001100110011001101",
    959 => "00111110010101111011100001100111",
    960 => "00111111011011011010000100000001",
    961 => "00111100011010000101111100001010",
    962 => "00111111010011101001010011100111",
    963 => "00111011000011011111111110010001",
    964 => "00111101110011001100110011001101",
    965 => "00111111011011011010000100000001",
    966 => "00111001110011100011101100011101",
    967 => "00111111000010110000000111000110",
    968 => "00111011011011010101111011011101",
    969 => "00111101110011001100110011001101",
    970 => "00111110011000010101100010101111",
    971 => "00111111011011011010000100000001",
    972 => "00111100011011000110110110100000",
    973 => "00111111010011011011101111010011",
    974 => "00111011000100010001101010100000",
    975 => "00111101110011001100110011001101",
    976 => "00111111011011011010000100000001",
    977 => "00111001110010100011100011100100",
    978 => "00111111000010100111011001011000",
    979 => "00111011011010011010110000010010",
    980 => "00111101110011001100110011001101",
    981 => "00111110011000101100100101000111",
    982 => "00111111011011011010000100000001",
    983 => "00111100011011010000110000000011",
    984 => "00111111010011011001101011110111",
    985 => "00111011000100011001010000101011",
    986 => "00111101110011001100110011001101",
    987 => "00111111011011011010000100000001",
    988 => "00111001110010011010010001000111",
    989 => "00111111000010100110000111111000",
    990 => "00111011011010010010001010100110",
    991 => "00111101110011001100110011001101",
    992 => "00111110011000101111111000111000",
    993 => "00111111011011011010000100000001",
    994 => "00111100011011010010001011011001",
    995 => "00111111010011011001011000111100",
    996 => "00111011000100011010010110110010",
    997 => "00111110011100111010000001111010",
    998 => "00111111100000000000000000000000",
    999 => "00111111101011100000011100001010");

  constant ans_lut : lut := (
    0 => "01000011000000000000000000000000",
    1 => "00000000000000000000000000000000",
    2 => "00111111011100001000111111111101",
    3 => "00111110101100101011011111111111",
    4 => "00111110101011110001110010010000",
    5 => "00111111010111011011010111111010",
    6 => "00111111000001100000100111111111",
    7 => "00111110111111111111111101000111",
    8 => "00111111010001000010010101001010",
    9 => "00111111010111110110010111111110",
    10 => "00111111001001001000111101111010",
    11 => "00111111010111110110010111111110",
    12 => "00111111010001000010010101001010",
    13 => "00111111010111110110010111111110",
    14 => "00111111001001001000111101111010",
    15 => "00000000000000000000000000000000",
    16 => "01000000000100000000000000000000",
    17 => "01000000010100000000000000000000",
    18 => "00000000000000000000000000000000",
    19 => "00111111100000000000000000000001",
    20 => "00000000000000000000000000000000",
    21 => "10111101110011001100110011001101",
    22 => "00000000000000000000000000000000",
    23 => "00111101110011001100110011001101",
    24 => "00111110110101100101110110110100",
    25 => "10111110000001011010100011011000",
    26 => "10111110000001100000101011000010",
    27 => "00111111011111011100111101010011",
    28 => "00111101110100000101100110000111",
    29 => "00111101110100000101100110000111",
    30 => "00111110110101101000100000000010",
    31 => "00111111011010111001100001111101",
    32 => "00111111100101011001101111100110",
    33 => "00111110110010000101000001010010",
    34 => "00111111001010011011001111001110",
    35 => "00111111010000000110110110010110",
    36 => "10111101101110011011111111101000",
    37 => "10111101101110100000000101011000",
    38 => "00111111011111101111000111100100",
    39 => "00111101110110000000111110000011",
    40 => "00111101110110000000111110000011",
    41 => "00111110110101110011011000100010",
    42 => "00111111011010011100101111001100",
    43 => "00111111100100110101101011101010",
    44 => "00111110110100001001010000111111",
    45 => "00111111001000010101010000110100",
    46 => "00111111001111101001101100011010",
    47 => "10111101101111001011111011010001",
    48 => "10111101101111010000001101111011",
    49 => "00111111011111101110100100010110",
    50 => "00111101110101111101101100100101",
    51 => "00111101110101111101101100100101",
    52 => "00111110110101110011000000110010",
    53 => "00111111011010011101011100101011",
    54 => "00111111100100110110100011100001",
    55 => "00111110110100000110000100111010",
    56 => "00111111001000011000001011111000",
    57 => "00111111001111101010010110110011",
    58 => "10111101101111001010110111000001",
    59 => "10111101101111001111001001011001",
    60 => "00111111011111101110100101001000",
    61 => "00111101110101111101110001010101",
    62 => "00111101110101111101110001010101",
    63 => "00111110110101110011000001011000",
    64 => "00111111011010011101011011101011",
    65 => "00111111100100110110100010010010",
    66 => "00111110110100000110001001011010",
    67 => "00111111001000011000000111110000",
    68 => "00111111001111101010010101111000",
    69 => "10111101101111001010111000100011",
    70 => "10111101101111001111001010111011",
    71 => "00111111011111101110100101001000",
    72 => "00111101110101111101110001001110",
    73 => "00111101110101111101110001001110",
    74 => "00111110110101110011000001010110",
    75 => "00111111011010011101011011101011",
    76 => "00111111100100110110100010010011",
    77 => "00111110110100000110001001010111",
    78 => "00111111000010010100101001000111",
    79 => "00111111110001001010010100100100",
    80 => "00111111110001001010010100100100",
    81 => "00111111100111101010011100000000",
    82 => "00000000000000000000000000000000",
    83 => "00111101110011001100110011001101",
    84 => "00111110110101100101110110110100",
    85 => "00111111011011001000001111011110",
    86 => "00111111100101101100110000011010",
    87 => "00111110110000111110111001001101",
    88 => "00111111001011101101000001000010",
    89 => "00111111001011101101000001000010",
    90 => "00111111010000010111011111111001",
    91 => "00111111001110010110101000011001",
    92 => "00111111010011110100000110101101",
    93 => "00111111001100001001100000000110",
    94 => "00111111010110100010111111111100",
    95 => "00111111010010001001101101110110",
    96 => "00111111001011101001011010111000",
    97 => "00111111010000000001110011100001",
    98 => "00111111001110110100110001010000",
    99 => "00111111010101110100101100101100",
    100 => "00111111010101110100101100101100",
    101 => "00111111010010000011010100111001",
    102 => "00111111001011110100001001011100",
    103 => "00111111010000010000011111100000",
    104 => "00111111001110101010110000110110",
    105 => "00111111010101110111110011011100",
    106 => "00111111010010000011110000100110",
    107 => "00111111001011110011011011001101",
    108 => "00111111010000001111100000000101",
    109 => "00111111001110101011011100001000",
    110 => "00111111010101110111100110010010",
    111 => "00111111010101110111100110010010",
    112 => "00111111010010000011101110110001",
    113 => "00111111001011110011011110010001",
    114 => "00111111010000001111100100010011",
    115 => "00111111001110101011011001001111",
    116 => "00111111010101110111100111001100",
    117 => "00111111010010000011101110111001",
    118 => "00111111001011110011011110000011",
    119 => "00111111010000001111100100000000",
    120 => "00111111001110101011011001011100",
    121 => "00111111010101110111100111000110",
    122 => "00111111010101110111100111000110",
    123 => "00111111010010000011101110111000",
    124 => "00111111001011110011011110000110",
    125 => "00111111010000001111100100000011",
    126 => "00111111001110101011011001011010",
    127 => "00111111010101110111100111001100",
    128 => "00111111010010000011101110111001",
    129 => "00111111001011110011011110000011",
    130 => "00111111010000001111100100000000",
    131 => "00111111001110101011011001011100",
    132 => "00111111010101110111100111000110",
    133 => "00111111010101110111100111000110",
    134 => "00111111010010000011101110111000",
    135 => "00111111001011110011011110000110",
    136 => "00111111010000001111100100000011",
    137 => "00111111001110101011011001011010",
    138 => "00111111101111011110000000110000",
    139 => "01000000000111101111000000011000",
    140 => "01000000000111101111000000011000",
    141 => "00111111110010011011011010000000",
    142 => "00000000000000000000000000000000",
    143 => "00111111011001100110011001101000",
    144 => "10111110100110011001100110011000",
    145 => "00000000000000000000000000000000",
    146 => "00111101110011001100110011001101",
    147 => "00111110110101100101110110110100",
    148 => "10111110110000111110111101011111",
    149 => "10111110110010010001000000100010",
    150 => "00111111011011001000001110100101",
    151 => "00111101111011111111000001000101",
    152 => "00111101111011111111000001000101",
    153 => "00111110110110110101111100111000",
    154 => "00111111011001011010011110010110",
    155 => "00111111100011100111101001000101",
    156 => "00111110111000100011110111000100",
    157 => "00111111000101010011011010110100",
    158 => "00111111001110111010110010111100",
    159 => "10111110100011110100000010111110",
    160 => "10111110100100010011000011100110",
    161 => "00111111011101011100011010011010",
    162 => "00111110000110010001011110000011",
    163 => "00111110000110010001011110000011",
    164 => "00111110111011100000001010110110",
    165 => "00111111011000000110001111101011",
    166 => "00111111100010001100011000101111",
    167 => "00111110111101100111100111100001",
    168 => "00111111000110000111101011000010",
    169 => "00111111001111001000000010011011",
    170 => "10111110100011100101100001111111",
    171 => "10111110100100000011111100001111",
    172 => "00111111011101011110100001010100",
    173 => "00111110000110010111111000010110",
    174 => "00111110000110010111111000010110",
    175 => "00111110111011100100000111100111",
    176 => "00111111011000000101101010110000",
    177 => "00111111100010001011110010011000",
    178 => "00111110111101101001101110000000",
    179 => "00111111000110001010001010101100",
    180 => "00111111001111001000101010001001",
    181 => "10111110100011100100110110000000",
    182 => "10111110100100000011001110011011",
    183 => "00111111011101011110100111101011",
    184 => "00111110000110011000001011100110",
    185 => "00111110000110011000001011100110",
    186 => "00111110111011100100010011100000",
    187 => "00111111011000000101101001000001",
    188 => "00111111100010001011110000100101",
    189 => "00111110111101101001110100010011",
    190 => "00111111000110001010010010001100",
    191 => "00111111001111001000101100000000",
    192 => "10111110100011100100110011111100",
    193 => "10111110100100000011001100010011",
    194 => "00111111011101011110100111111110",
    195 => "00111110000110011000001100100000",
    196 => "00111110000110011000001100100000",
    197 => "00111110111011100100010100000001",
    198 => "00111111011000000101101000111100",
    199 => "00111111100010001011110000100000",
    200 => "00111110111101101001110100100100",
    201 => "00111111000010111101001000111000",
    202 => "00111111110001011110100100011100",
    203 => "00111111110001011110100100011100",
    204 => "00111111100111110010100101111011",
    205 => "00111111001100110011001100110100",
    206 => "00000000000000000000000000000000",
    207 => "00111101110011001100110011001101",
    208 => "00111110110101100101110110110100",
    209 => "00111111010010110010000001111101",
    210 => "00111111011010101001001011010101",
    211 => "00111111000110111101100000101010",
    212 => "00111110100010100010100011110001",
    213 => "00111110100010100010100011110001",
    214 => "00111111000101110001011110110110",
    215 => "00111111010110001010110001101100",
    216 => "00111111100000010010100101000010",
    217 => "00111111000010000101101110111110",
    218 => "00111111010010000000000110010000",
    219 => "00111111010001011110111101110011",
    220 => "00111111000100001110111110100100",
    221 => "00111111000110100001000101111000",
    222 => "00111111010100110000100110110010",
    223 => "00111110111011111110010110110110",
    224 => "00111110111011111110010110110110",
    225 => "00111111001100101011000010111110",
    226 => "00111111010010010011110100110100",
    227 => "00111111011001110111110111000110",
    228 => "00111111000111100100011101011010",
    229 => "00111111010110110111001001011010",
    230 => "00111111010010001100011100111010",
    231 => "00111111000011001101001100010110",
    232 => "00111111000101010001110100000001",
    233 => "00111111010101011100110011101001",
    234 => "00111110111100011010001010100000",
    235 => "00111110111100011010001010100000",
    236 => "00111111001100110000000110010010",
    237 => "00111111010010001111100010111100",
    238 => "00111111011001110000111011110101",
    239 => "00111111000111101001111001101000",
    240 => "00111111010110110111111101011100",
    241 => "00111111010010001100100011111100",
    242 => "00111111000011001101000001101110",
    243 => "00111111000101010001100111010100",
    244 => "00111111010101011100111010101000",
    245 => "00111110111100011010001110011000",
    246 => "00111110111100011010001110011000",
    247 => "00111111001100110000000111000000",
    248 => "00111111010010001111100010011000",
    249 => "00111111011001110000111010111010",
    250 => "00111111000111101001111010010110",
    251 => "00111111010110110111111101101100",
    252 => "00111111010010001100100011111110",
    253 => "00111111000011001101000001101100",
    254 => "00111111000101010001100111010001",
    255 => "00111111010101011100111010101010",
    256 => "00111110111100011010001110100101",
    257 => "00111110111100011010001110100101",
    258 => "00111111001100110000000111000011",
    259 => "00111111010010001111100010010101",
    260 => "00111111011001110000111010110110",
    261 => "00111111000111101001111010011001",
    262 => "00111111100100001000111100000011",
    263 => "01000000000010000100011110000010",
    264 => "01000000000010000100011110000010",
    265 => "00111111101110101100100000101111",
    266 => "00000000000000000000000000000000",
    267 => "00111101110011001100110011001101",
    268 => "00111110110101100101110110110100",
    269 => "10111111000110111101100010100001",
    270 => "10111111001001111000110101110001",
    271 => "00111111010010110010000000100010",
    272 => "00111110001000101011000101101010",
    273 => "00111110001000101011000101101010",
    274 => "00111110111100111110111001111010",
    275 => "00111111010111111001110000010100",
    276 => "00111111100001111111011110101111",
    277 => "00111110111110010100110010100010",
    278 => "00111111000111000111101111111000",
    279 => "00111111001111010111101001111110",
    280 => "10111110111001011111101011110010",
    281 => "10111110111011101000001101110000",
    282 => "00111111011001001011100110000010",
    283 => "00111110100000100100111001000101",
    284 => "00111110100000100100111001000101",
    285 => "00111111000100111101100010100110",
    286 => "00111111010110011011100011010111",
    287 => "00111111100000100010011100000000",
    288 => "00111111000001101010110100101100",
    289 => "00111111010000111101110011011100",
    290 => "00111111010001010100010010001000",
    291 => "10111110110101101101010000000110",
    292 => "10111110110111011011000010111100",
    293 => "00111111011010000110000010100101",
    294 => "00111110100001101110011001010010",
    295 => "00111110100001101110011001010010",
    296 => "00111111000101011100010111001001",
    297 => "00111111010110010001110100110010",
    298 => "00111111100000011001001101111011",
    299 => "00111111000001111010011111000000",
    300 => "00111111010001100101110001110110",
    301 => "00111111010001011010110001010010",
    302 => "10111110110101011111001111011110",
    303 => "10111110110111001011100111100110",
    304 => "00111111011010001001010001001111",
    305 => "00111110100001110010000111000011",
    306 => "00111110100001110010000111000011",
    307 => "00111111000101011101111000101110",
    308 => "00111111010110010001010100111010",
    309 => "00111111100000011000101111110101",
    310 => "00111111000001111011010010000010",
    311 => "00111111010001100111101101100010",
    312 => "00111111010001011011000101001010",
    313 => "10111110110101011110100100010100",
    314 => "10111110110111001010111000000110",
    315 => "00111111011010001001011011001010",
    316 => "00111110100001110010010010010110",
    317 => "00111110100001110010010010010110",
    318 => "00111111000101011101111101010111",
    319 => "00111111010110010001010011011001",
    320 => "00111111100000011000101110011010",
    321 => "00111111000001111011010100011100",
    322 => "00111111010101101101101111110011",
    323 => "00111111111010110110110111111010",
    324 => "00111111111010110110110111111010",
    325 => "00111111101011011001100000100101",
    326 => "00111111000000000000000000000000",
    327 => "00000000000000000000000000000000",
    328 => "00111101110011001100110011001101",
    329 => "00111110110101100101110110110100",
    330 => "00111111000110111101100010100011",
    331 => "00111111001001111000110101110100",
    332 => "00111111010010110010000000100000",
    333 => "00111110001000101011000101101100",
    334 => "00111110001000101011000101101100",
    335 => "00111110111100111110111001111010",
    336 => "00111111010111111001110000010100",
    337 => "00111111100001111111011110101111",
    338 => "00111110111110010100110010100010",
    339 => "00111111000111000111101111111010",
    340 => "00111111001111010111101001111110",
    341 => "00111110111001011111101011110101",
    342 => "00111110111011101000001101110011",
    343 => "00111111011001001011100110000001",
    344 => "00111110100000100100111001001001",
    345 => "00111110100000100100111001001001",
    346 => "00111111000100111101100010101000",
    347 => "00111111010110011011100011010110",
    348 => "00111111100000100010011011111111",
    349 => "00111111000001101010110100101110",
    350 => "00111111010000111101110011011100",
    351 => "00111111010001010100010010001000",
    352 => "00111110110101101101010000001001",
    353 => "00111110110111011011000010111111",
    354 => "00111111011010000110000010100101",
    355 => "00111110100001101110011001010011",
    356 => "00111110100001101110011001010011",
    357 => "00111111000101011100010111001011",
    358 => "00111111010110010001110100110010",
    359 => "00111111100000011001001101111100",
    360 => "00111111000001111010011110111110",
    361 => "00111111010001100101110001111110",
    362 => "00111111010001011010110001010011",
    363 => "00111110110101011111001111100000",
    364 => "00111110110111001011100111100111",
    365 => "00111111011010001001010001001110",
    366 => "00111110100001110010000111001001",
    367 => "00111110100001110010000111001001",
    368 => "00111111000101011101111000110000",
    369 => "00111111010110010001010100111000",
    370 => "00111111100000011000101111110100",
    371 => "00111111000001111011010010000011",
    372 => "00111111010001100111101101100100",
    373 => "00111111010001011011000101001010",
    374 => "00111110110101011110100100010111",
    375 => "00111110110111001010111000001001",
    376 => "00111111011010001001011011001001",
    377 => "00111110100001110010010010011001",
    378 => "00111110100001110010010010011001",
    379 => "00111111000101011101111101011010",
    380 => "00111111010110010001010011011001",
    381 => "00111111100000011000101110011010",
    382 => "00111111000001111011010100011100",
    383 => "00111111010101101101101111111010",
    384 => "00111111111010110110110111111101",
    385 => "00111111111010110110110111111101",
    386 => "00111111101011011001100000100110",
    387 => "00000000000000000000000000000000",
    388 => "00111111011001100110011001101000",
    389 => "10111111001100110011001100110010",
    390 => "00000000000000000000000000000000",
    391 => "00111101110011001100110011001101",
    392 => "00111110110101100101110110110100",
    393 => "10111111010010110010000001011000",
    394 => "10111111011010101001001011010011",
    395 => "00111111000111000000110001111010",
    396 => "00111110100010100010100100010100",
    397 => "00111110100010100010100100010100",
    398 => "00111111000101110001011111000101",
    399 => "00111111010110001010110001101000",
    400 => "00111111100000010010100100111110",
    401 => "00111111000010000101101111000101",
    402 => "00111111010010000000000110100100",
    403 => "00111111010001011110111101110111",
    404 => "10111111000100001110111110100000",
    405 => "10111111000110100001000101110010",
    406 => "00111111010100110000100110110100",
    407 => "00111110111011111110010110111101",
    408 => "00111110111011111110010110111101",
    409 => "00111111001100101011000011000000",
    410 => "00111111010010010011110100110010",
    411 => "00111111011001110111110111000100",
    412 => "00111111000111100100011101011011",
    413 => "00111111010110110111001001011010",
    414 => "00111111010010001100011100111010",
    415 => "10111111000011001101001100010100",
    416 => "10111111000101010001110011111111",
    417 => "00111111010101011100110011101011",
    418 => "00111110111100011010001010010110",
    419 => "00111110111100011010001010010110",
    420 => "00111111001100110000000110010001",
    421 => "00111111010010001111100010111111",
    422 => "00111111011001110000111011111001",
    423 => "00111111000111101001111001100100",
    424 => "00111111010110110111111101100010",
    425 => "00111111010010001100100011111100",
    426 => "10111111000011001101000001101110",
    427 => "10111111000101010001100111010010",
    428 => "00111111010101011100111010101001",
    429 => "00111110111100011010001110011101",
    430 => "00111110111100011010001110011101",
    431 => "00111111001100110000000111000000",
    432 => "00111111010010001111100010010101",
    433 => "00111111011001110000111010110110",
    434 => "00111111000111101001111010011001",
    435 => "00111111010110110111111101100010",
    436 => "00111111010010001100100011111100",
    437 => "10111111000011001101000001101110",
    438 => "10111111000101010001100111010010",
    439 => "00111111010101011100111010101001",
    440 => "00111110111100011010001110011101",
    441 => "00111110111100011010001110011101",
    442 => "00111111001100110000000111000000",
    443 => "00111111010010001111100010010101",
    444 => "00111111011001110000111010110110",
    445 => "00111111000111101001111010011001",
    446 => "00111111100100001000111011111110",
    447 => "01000000000010000100011101111111",
    448 => "01000000000010000100011101111111",
    449 => "00111111101110101100100000101101",
    450 => "00111110100110011001100110011010",
    451 => "00000000000000000000000000000000",
    452 => "00111101110011001100110011001101",
    453 => "00111110110101100101110110110100",
    454 => "00111110110000111110111101100001",
    455 => "00111110110010010001000000100100",
    456 => "00111111011011001000001110100101",
    457 => "00111101111011111111000001000110",
    458 => "00111101111011111111000001000110",
    459 => "00111110110110110101111100111000",
    460 => "00111111011001011010011110010110",
    461 => "00111111100011100111101001000101",
    462 => "00111110111000100011110111000100",
    463 => "00111111000101010011011010110101",
    464 => "00111111001110111010110010111100",
    465 => "00111110100011110100000011000000",
    466 => "00111110100100010011000011101000",
    467 => "00111111011101011100011010011010",
    468 => "00111110000110010001011110000100",
    469 => "00111110000110010001011110000100",
    470 => "00111110111011100000001010111001",
    471 => "00111111011000000110001111101011",
    472 => "00111111100010001100011000101111",
    473 => "00111110111101100111100111100001",
    474 => "00111111000110000111101011000011",
    475 => "00111111001111001000000010011011",
    476 => "00111110100011100101100010000001",
    477 => "00111110100100000011111100010001",
    478 => "00111111011101011110100001010100",
    479 => "00111110000110010111111000011000",
    480 => "00111110000110010111111000011000",
    481 => "00111110111011100100000111101010",
    482 => "00111111011000000101101010110000",
    483 => "00111111100010001011110010011000",
    484 => "00111110111101101001101110000000",
    485 => "00111111000110001010001010101110",
    486 => "00111111001111001000101010001001",
    487 => "00111110100011100100110110000010",
    488 => "00111110100100000011001110011101",
    489 => "00111111011101011110100111101011",
    490 => "00111110000110011000001011101000",
    491 => "00111110000110011000001011101000",
    492 => "00111110111011100100010011100000",
    493 => "00111111011000000101101001000001",
    494 => "00111111100010001011110000100101",
    495 => "00111110111101101001110100010011",
    496 => "00111111000110001010010010001110",
    497 => "00111111001111001000101100000000",
    498 => "00111110100011100100110011111110",
    499 => "00111110100100000011001100010101",
    500 => "00111111011101011110100111111110",
    501 => "00111110000110011000001100100010",
    502 => "00111110000110011000001100100010",
    503 => "00111110111011100100010100000100",
    504 => "00111111011000000101101000111100",
    505 => "00111111100010001011110000011111",
    506 => "00111110111101101001110100100111",
    507 => "00111111000010111101001000111011",
    508 => "00111111110001011110100100011110",
    509 => "00111111110001011110100100011110",
    510 => "00111111100111110010100101111011",
    511 => "00000000000000000000000000000000",
    512 => "00111101110011001100110011001101",
    513 => "00111110110101100101110110110100",
    514 => "10111111011011001010101110011111",
    515 => "10111111100101101100110000011010",
    516 => "00111110110001011100100001110101",
    517 => "00111111001011101101100011000110",
    518 => "00111111001011101101100011000110",
    519 => "00111111010000010111100110101001",
    520 => "00111111001110010110011111011000",
    521 => "00111111010011110011111001100101",
    522 => "00111111001100001001101001100111",
    523 => "00111111010110100010111101110110",
    524 => "00111111010010001001101101100100",
    525 => "10111111001011101001011011010110",
    526 => "10111111010000000001110100001010",
    527 => "00111111001110110100110000110011",
    528 => "00111111010101110100101100110000",
    529 => "00111111010101110100101100110000",
    530 => "00111111010010000011010100111010",
    531 => "00111111001011110100001001011011",
    532 => "00111111010000010000011111011110",
    533 => "00111111001110101010110000111000",
    534 => "00111111010101110111110011011000",
    535 => "00111111010010000011110000100110",
    536 => "10111111001011110011011011001101",
    537 => "10111111010000001111100000000101",
    538 => "00111111001110101011011100001000",
    539 => "00111111010101110111100110001110",
    540 => "00111111010101110111100110001110",
    541 => "00111111010010000011101110110000",
    542 => "00111111001011110011011110010011",
    543 => "00111111010000001111100100010101",
    544 => "00111111001110101011011001001101",
    545 => "00111111010101110111100111010100",
    546 => "00111111010010000011101110111010",
    547 => "10111111001011110011011101111111",
    548 => "10111111010000001111100011111010",
    549 => "00111111001110101011011001100000",
    550 => "00111111010101110111100110111100",
    551 => "00111111010101110111100110111100",
    552 => "00111111010010000011101110110111",
    553 => "00111111001011110011011110000111",
    554 => "00111111010000001111100100000101",
    555 => "00111111001110101011011001011001",
    556 => "00111111010101110111100111000110",
    557 => "00111111010010000011101110111000",
    558 => "10111111001011110011011110000100",
    559 => "10111111010000001111100100000001",
    560 => "00111111001110101011011001011100",
    561 => "00111111010101110111100111000100",
    562 => "00111111010101110111100111000100",
    563 => "00111111010010000011101110111000",
    564 => "00111111001011110011011110000110",
    565 => "00111111010000001111100100000011",
    566 => "00111111001110101011011001011010",
    567 => "00111111101111011110000000101110",
    568 => "01000000000111101111000000010111",
    569 => "01000000000111101111000000010111",
    570 => "00111111110010011011011001111111",
    571 => "00111101110011001100110011001101",
    572 => "00000000000000000000000000000000",
    573 => "00111101110011001100110011001101",
    574 => "00111110110101100101110110110100",
    575 => "00111110000001011010100011011000",
    576 => "00111110000001100000101011000010",
    577 => "00111111011111011100111101010011",
    578 => "00111101110100000101100110000111",
    579 => "00111101110100000101100110000111",
    580 => "00111110110101101000100000000010",
    581 => "00111111011010111001100001111101",
    582 => "00111111100101011001101111100110",
    583 => "00111110110010000101000001010010",
    584 => "00111111001010011011001111001110",
    585 => "00111111010000000110110110010110",
    586 => "00111101101110011011111111101000",
    587 => "00111101101110100000000101011000",
    588 => "00111111011111101111000111100100",
    589 => "00111101110110000000111110000011",
    590 => "00111101110110000000111110000011",
    591 => "00111110110101110011011000100010",
    592 => "00111111011010011100101111001100",
    593 => "00111111100100110101101011101010",
    594 => "00111110110100001001010000111111",
    595 => "00111111001000010101010000110100",
    596 => "00111111001111101001101100011010",
    597 => "00111101101111001011111011010001",
    598 => "00111101101111010000001101111011",
    599 => "00111111011111101110100100010110",
    600 => "00111101110101111101101100100101",
    601 => "00111101110101111101101100100101",
    602 => "00111110110101110011000000110010",
    603 => "00111111011010011101011100101011",
    604 => "00111111100100110110100011100001",
    605 => "00111110110100000110000100111010",
    606 => "00111111001000011000001011111000",
    607 => "00111111001111101010010110110011",
    608 => "00111101101111001010110111000001",
    609 => "00111101101111001111001001011001",
    610 => "00111111011111101110100101001000",
    611 => "00111101110101111101110001010101",
    612 => "00111101110101111101110001010101",
    613 => "00111110110101110011000001011000",
    614 => "00111111011010011101011011101011",
    615 => "00111111100100110110100010010010",
    616 => "00111110110100000110001001011010",
    617 => "00111111001000011000000111110000",
    618 => "00111111001111101010010101111000",
    619 => "00111101101111001010111000100011",
    620 => "00111101101111001111001010111011",
    621 => "00111111011111101110100101001000",
    622 => "00111101110101111101110001001110",
    623 => "00111101110101111101110001001110",
    624 => "00111110110101110011000001010110",
    625 => "00111111011010011101011011101011",
    626 => "00111111100100110110100010010011",
    627 => "00111110110100000110001001010111",
    628 => "00111111000010010100101001000111",
    629 => "00111111110001001010010100100100",
    630 => "00111111110001001010010100100100",
    631 => "00111111100111101010011100000000",
    632 => "00000000000000000000000000000000",
    633 => "00111111001100110011001100110110",
    634 => "10111101110011001100110011000000",
    635 => "00000000000000000000000000000000",
    636 => "00111101110011001100110011001101",
    637 => "00111110110101100101110110110100",
    638 => "10111110000001011010100011010000",
    639 => "10111110000001100000101010111010",
    640 => "00111111011111011100111101010011",
    641 => "00111101110100000101100110000110",
    642 => "00111101110100000101100110000110",
    643 => "00111110110101101000100000000010",
    644 => "00111111010010011111111110001100",
    645 => "00111111011010001011100110100000",
    646 => "00111111000111010100111010011000",
    647 => "00111110100010010001000011100000",
    648 => "00111111000101101010011101101010",
    649 => "10111101111001010110001010111110",
    650 => "10111101111001011101111000111000",
    651 => "00111111011111100110001110100001",
    652 => "00111101110100111100001111110001",
    653 => "00111101110100111100001111110001",
    654 => "00111110110101101100100000011100",
    655 => "00111111010010001111110111110100",
    656 => "00111111011001110001011101100100",
    657 => "00111111000111101001011111001000",
    658 => "00111110100010000011010110011001",
    659 => "00111111000101100100111010110111",
    660 => "10111101111001011001010000010010",
    661 => "10111101111001100000111111011101",
    662 => "00111111011111100110001011101110",
    663 => "00111101110100111011101111010000",
    664 => "00111101110100111011101111010000",
    665 => "00111110110101101100011101101100",
    666 => "00111111010010010000000001000011",
    667 => "00111111011001110001101100100000",
    668 => "00111111000111101001010011011010",
    669 => "00111110100010000011011101101111",
    670 => "00111111000101100100111101111000",
    671 => "10111101111001011001001110101001",
    672 => "10111101111001100000111101110011",
    673 => "00111111011111100110001011101111",
    674 => "00111101110100111011101111100010",
    675 => "00111101110100111011101111100010",
    676 => "00111110110101101100011101101110",
    677 => "00111111010010010000000000111110",
    678 => "00111111011001110001101100011001",
    679 => "00111111000111101001010011100000",
    680 => "00111110100010000011011101101100",
    681 => "00111111000101100100111101110101",
    682 => "10111101111001011001001110101001",
    683 => "10111101111001100000111101110011",
    684 => "00111111011111100110001011101111",
    685 => "00111101110100111011101111100010",
    686 => "00111101110100111011101111100010",
    687 => "00111110110101101100011101101110",
    688 => "00111111010010010000000000111110",
    689 => "00111111011001110001101100011001",
    690 => "00111111000111101001010011100000",
    691 => "00111110001011010111111111111100",
    692 => "00111111100101011011000000000000",
    693 => "00111111100101011011000000000000",
    694 => "00111111100010100110101101101110",
    695 => "00111111011001100110011001101000",
    696 => "00000000000000000000000000000000",
    697 => "00111101110011001100110011001101",
    698 => "00111110110101100101110110110100",
    699 => "00111111011011001000001111011110",
    700 => "00111111100101101100110000011011",
    701 => "00111110110000111110111001001001",
    702 => "00111111001011101101000001001000",
    703 => "00111111001011101101000001001000",
    704 => "00111111010000010111011111111011",
    705 => "00111111000101101100001000001010",
    706 => "00111111001000010011001100010100",
    707 => "00111111010011101110110010100010",
    708 => "00111110111011001101000111000001",
    709 => "00111111001100100001111101011000",
    710 => "00111111010010011011011010101010",
    711 => "00111111011010000100001011110011",
    712 => "00111111000111011010110000101100",
    713 => "00111111010110110101100001111000",
    714 => "00111111010110110101100001111000",
    715 => "00111111010010001100001110111011",
    716 => "00111111000011001101100001011001",
    717 => "00111111000101010010001101001111",
    718 => "00111111010101011100100101110010",
    719 => "00111110111100011010000010001101",
    720 => "00111111001100110000000100110011",
    721 => "00111111010010001111100100001111",
    722 => "00111111011001110000111101111011",
    723 => "00111111000111101001110111111110",
    724 => "00111111010110110111111101010110",
    725 => "00111111010110110111111101010110",
    726 => "00111111010010001100100011111011",
    727 => "00111111000011001101000001110010",
    728 => "00111111000101010001100111010111",
    729 => "00111111010101011100111010100110",
    730 => "00111110111100011010001110100101",
    731 => "00111111001100110000000111000011",
    732 => "00111111010010001111100010010101",
    733 => "00111111011001110000111010110110",
    734 => "00111111000111101001111010011001",
    735 => "00111111010110110111111101100110",
    736 => "00111111010110110111111101100110",
    737 => "00111111010010001100100011111101",
    738 => "00111111000011001101000001101110",
    739 => "00111111000101010001100111010100",
    740 => "00111111010101011100111010101000",
    741 => "00111110111100011010001110100010",
    742 => "00111111001100110000000111000010",
    743 => "00111111010010001111100010010101",
    744 => "00111111011001110000111010110110",
    745 => "00111111000111101001111010011001",
    746 => "00111111010110110111111101100100",
    747 => "00111111010110110111111101100100",
    748 => "00111111010010001100100011111101",
    749 => "00111111000011001101000001101110",
    750 => "00111111000101010001100111010100",
    751 => "00111111010101011100111010101000",
    752 => "00111111100100001000111100000001",
    753 => "01000000000010000100011110000000",
    754 => "01000000000010000100011110000000",
    755 => "00111111101110101100100000101110",
    756 => "00000000000000000000000000000000",
    757 => "00111101110011001100110011001101",
    758 => "00111110110101100101110110110100",
    759 => "10111110110000111110111101011111",
    760 => "10111110110010010001000000100010",
    761 => "00111111011011001000001110100101",
    762 => "00111101111011111111000001000101",
    763 => "00111101111011111111000001000101",
    764 => "00111110110110110101111100111000",
    765 => "00111111010000110000001000001010",
    766 => "00111111010111011010000111000100",
    767 => "00111111001001011110100011111000",
    768 => "00111110100001100000100111000111",
    769 => "00111111000101010110101011010111",
    770 => "10111110101010011010010100011111",
    771 => "10111110101011001110100111001001",
    772 => "00111111011100011000101000100101",
    773 => "00111110000001110111010111010001",
    774 => "00111110000001110111010111010001",
    775 => "00111110111000110110101101111010",
    776 => "00111111001111110110110100110000",
    777 => "00111111010110000010100100101010",
    778 => "00111111001010100000101000011110",
    779 => "00111110100010001111111110100000",
    780 => "00111111000101101010000001110100",
    781 => "10111110101010010010110000110000",
    782 => "10111110101011000110100110100010",
    783 => "00111111011100011001111101011000",
    784 => "00111110000001111111101010111100",
    785 => "00111110000001111111101010111100",
    786 => "00111110111000111011011111011010",
    787 => "00111111001111110101011011011000",
    788 => "00111111010110000000011101110100",
    789 => "00111111001010100010001101010010",
    790 => "00111110100010010010011000101010",
    791 => "00111111000101101010111111111100",
    792 => "10111110101010010010011000000010",
    793 => "10111110101011000110001100010101",
    794 => "00111111011100011010000001101110",
    795 => "00111110000010000000000101101100",
    796 => "00111110000010000000000101101100",
    797 => "00111110111000111011101110110011",
    798 => "00111111001111110101010110111101",
    799 => "00111111010110000000010111001000",
    800 => "00111111001010100010010010010010",
    801 => "00111110100010010010100000100011",
    802 => "00111111000101101011000011001000",
    803 => "10111110101010010010010110110001",
    804 => "10111110101011000110001011000000",
    805 => "00111111011100011010000001111100",
    806 => "00111110000010000000000111000100",
    807 => "00111110000010000000000111000100",
    808 => "00111110111000111011101111100111",
    809 => "00111111001111110101010110101101",
    810 => "00111111010110000000010110110001",
    811 => "00111111001010100010010010100011",
    812 => "00111110010011011000010101110000",
    813 => "00111111100110011011000010101110",
    814 => "00111111100110011011000010101110",
    815 => "00111111100011000100001000010100",
    816 => "00111111001100110011001100110100",
    817 => "00000000000000000000000000000000",
    818 => "00111101110011001100110011001101",
    819 => "00111110110101100101110110110100",
    820 => "00111111010010110010000001111101",
    821 => "00111111011010101001001011010101",
    822 => "00111111000110111101100000101010",
    823 => "00111110100010100010100011110001",
    824 => "00111110100010100010100011110001",
    825 => "00111111000101110001011110110110",
    826 => "00111111001101001110110100100000",
    827 => "00111111010010001110101011011011",
    828 => "00111111001101010011010000010100",
    829 => "00111110101111010000110001011100",
    830 => "00111111001001111001001000011001",
    831 => "00111111001011010100101111111111",
    832 => "00111111001111100101101001001001",
    833 => "00111111001111000111110110011010",
    834 => "00111110110100110001011010010000",
    835 => "00111110110100110001011010010000",
    836 => "00111111001011001110001010010011",
    837 => "00111111001010011110100100101110",
    838 => "00111111001110011100101001111100",
    839 => "00111111001111111000101001011010",
    840 => "00111110110110010110001001101001",
    841 => "00111111001011100100000011101100",
    842 => "00111111001010001111001110010101",
    843 => "00111111001110001000001011110110",
    844 => "00111111010000000110001010010110",
    845 => "00111110110110101110110110010010",
    846 => "00111110110110101110110110010010",
    847 => "00111111001011101001010001111010",
    848 => "00111111001010001011011110010110",
    849 => "00111111001110000011001100101011",
    850 => "00111111010000001001011100010100",
    851 => "00111110110110110100101010010011",
    852 => "00111111001011101010100000000010",
    853 => "00111111001010001010100101111001",
    854 => "00111111001110000010000001101001",
    855 => "00111111010000001010001101101000",
    856 => "00111110110110110110000001000011",
    857 => "00111110110110110110000001000011",
    858 => "00111111001011101010110010010000",
    859 => "00111111001010001010011000110000",
    860 => "00111111001110000001110000001011",
    861 => "00111111010000001010011001000111",
    862 => "00111110110110110110010101001101",
    863 => "00111111001011101010110110011110",
    864 => "00111111001010001010010101101010",
    865 => "00111111001110000001101100000101",
    866 => "00111111010000001010011011110011",
    867 => "00111110110110110110011001110101",
    868 => "00111110110110110110011001110101",
    869 => "00111111001011101010110111011100",
    870 => "00111111001010001010010100111111",
    871 => "00111111001110000001101011001011",
    872 => "00111111010000001010011100011010",
    873 => "00111111001010000011001101100110",
    874 => "00111111110101000001100110110011",
    875 => "00111111110101000001100110110011",
    876 => "00111111101001001100010011100010",
    877 => "00000000000000000000000000000000",
    878 => "00111111001100110011001100110110",
    879 => "10111110111111111111111111111110",
    880 => "00000000000000000000000000000000",
    881 => "00111101110011001100110011001101",
    882 => "00111110110101100101110110110100",
    883 => "10111111000110111101100010100001",
    884 => "10111111001001111000110101110001",
    885 => "00111111010010110010000000100010",
    886 => "00111110001000101011000101101010",
    887 => "00111110001000101011000101101010",
    888 => "00111110111100111110111001111010",
    889 => "00111111001111000100111110011010",
    890 => "00111111010100111000000101001100",
    891 => "00111111001011010111111000011111",
    892 => "00111110100100101111101101100110",
    893 => "00111111000110100111101011011001",
    894 => "10111111000001110000100100001100",
    895 => "10111111000011100011110111000101",
    896 => "00111111010110010111111111110100",
    897 => "00111110010101111011100001011110",
    898 => "00111110010101111011100001011110",
    899 => "00111111000010010011011011100101",
    900 => "00111111001110001111001100100001",
    901 => "00111111010011101001010011101010",
    902 => "00111111001100010001010100000000",
    903 => "00111110101010001100011101101001",
    904 => "00111111001000011101001100010000",
    905 => "10111111000001000100011011010100",
    906 => "10111111000010110000000111000100",
    907 => "00111111010110110010111111101001",
    908 => "00111110011000010101100010101110",
    909 => "00111110011000010101100010101110",
    910 => "00111111000010111010110010011000",
    911 => "00111111001110000101110100101110",
    912 => "00111111010011011011101111010011",
    913 => "00111111001100011011000110010110",
    914 => "00111110101011000110100001011111",
    915 => "00111111001000101110110000110011",
    916 => "10111111000000111100111101100000",
    917 => "10111111000010100111011001010110",
    918 => "00111111010110110111011111000110",
    919 => "00111110011000101100100101000111",
    920 => "00111110011000101100100101000111",
    921 => "00111111000011000000100010010000",
    922 => "00111111001110000100011001110000",
    923 => "00111111010011011001101011110111",
    924 => "00111111001100011100100100111111",
    925 => "00111110101011001111000000001011",
    926 => "00111111001000110001010010010011",
    927 => "10111111000000111011110111101000",
    928 => "10111111000010100110000111110110",
    929 => "00111111010110111000001001000000",
    930 => "00111110011000101111111000110100",
    931 => "00111110011000101111111000110100",
    932 => "00111111000011000001010110111000",
    933 => "00111111001110000100001100101001",
    934 => "00111111010011011001011000111100",
    935 => "00111111001100011100110010100110",
    936 => "00111110101110000001110000100001",
    937 => "00111111101011100000011100001000",
    938 => "00111111101011100000011100001000",
    939 => "00111111100101010011111111110101",
    940 => "00111111000000000000000000000000",
    941 => "00000000000000000000000000000000",
    942 => "00111101110011001100110011001101",
    943 => "00111110110101100101110110110100",
    944 => "00111111000110111101100010100011",
    945 => "00111111001001111000110101110100",
    946 => "00111111010010110010000000100000",
    947 => "00111110001000101011000101101100",
    948 => "00111110001000101011000101101100",
    949 => "00111110111100111110111001111010",
    950 => "00111111001111000100111110011010",
    951 => "00111111010100111000000101001100",
    952 => "00111111001011010111111000011111",
    953 => "00111110100100101111101101100111",
    954 => "00111111000110100111101011011010",
    955 => "00111111000001110000100100001110",
    956 => "00111111000011100011110111000111",
    957 => "00111111010110010111111111110011",
    958 => "00111110010101111011100001100111",
    959 => "00111110010101111011100001100111",
    960 => "00111111000010010011011011100110",
    961 => "00111111001110001111001100011111",
    962 => "00111111010011101001010011100111",
    963 => "00111111001100010001010100000010",
    964 => "00111110101010001100011101101000",
    965 => "00111111001000011101001100001110",
    966 => "00111111000001000100011011010110",
    967 => "00111111000010110000000111000110",
    968 => "00111111010110110010111111101000",
    969 => "00111110011000010101100010101111",
    970 => "00111110011000010101100010101111",
    971 => "00111111000010111010110010011000",
    972 => "00111111001110000101110100101110",
    973 => "00111111010011011011101111010011",
    974 => "00111111001100011011000110010110",
    975 => "00111110101011000110100001011111",
    976 => "00111111001000101110110000110011",
    977 => "00111111000000111100111101100001",
    978 => "00111111000010100111011001011000",
    979 => "00111111010110110111011111000101",
    980 => "00111110011000101100100101000111",
    981 => "00111110011000101100100101000111",
    982 => "00111111000011000000100010010000",
    983 => "00111111001110000100011001110000",
    984 => "00111111010011011001101011110111",
    985 => "00111111001100011100100100111111",
    986 => "00111110101011001111000000001011",
    987 => "00111111001000110001010010010011",
    988 => "00111111000000111011110111101010",
    989 => "00111111000010100110000111111000",
    990 => "00111111010110111000001001000000",
    991 => "00111110011000101111111000111000",
    992 => "00111110011000101111111000111000",
    993 => "00111111000011000001010110111010",
    994 => "00111111001110000100001100101001",
    995 => "00111111010011011001011000111100",
    996 => "00111111001100011100110010100110",
    997 => "00111110101110000001110000100110",
    998 => "00111111101011100000011100001010",
    999 => "00111111101011100000011100001010");


  component fadd is
    port (A : in std_logic_vector (31 downto 0);
          B : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          C : out std_logic_vector (31 downto 0));
  end component fadd;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal s_b : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (3 downto 0) of std_logic_vector (31 downto 0);
  signal cc : buff := (others => (others => '0'));
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');

  signal i_isRunning : std_logic := 'U';
  signal i_result : std_logic := '1';
begin  -- architecture fadd_tb

  i_fadd : fadd port map (s_a,s_b,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk) is
    variable ss : character;
    variable count : integer := 4;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      case state is
        when "00" =>
          state <= "01";
        when "01" =>
          state <= "11";
        when "11" =>
          state <= "10";
        when others =>
          state <= "00";
      end case;
      s_a <= a_lut (addr);
      s_b <= b_lut (addr);
      cc(conv_integer(state)) <= ans_lut (addr);      
        ccc <= cc (conv_integer (state));
      if i_isRunning = '1' then  -- rising clock edge
        if (ccc = c or state /= "00") and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 5 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;
  end process ram_loop;

end architecture;
