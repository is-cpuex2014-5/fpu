library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity finv_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity finv_tb;

architecture testbench of finv_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "01110001110111100011010110101110",
    1 => "11111010101110001010000010101001",
    2 => "11001011110100010100001100010110",
    3 => "01101110000101110100110101100101",
    4 => "11100001000011011101010000111111",
    5 => "00110110100001010000100001100110",
    6 => "01010000100011110100111110011011",
    7 => "01000101100110011011110111001001",
    8 => "10011011010001100111100101110001",
    9 => "10001110000010101101101011111000",
    10 => "10100011011000000001110001011111",
    11 => "10111110110001001100000110111111",
    12 => "10110000100000101110111000001010",
    13 => "00101010110001100101001011111111",
    14 => "11001111000101100010000100110011",
    15 => "01111011100000110001111010100011",
    16 => "01101000110101011101110001101100",
    17 => "00001001000010100011101110011110",
    18 => "01000001111110111011001101111001",
    19 => "01111010100100101100010101011001",
    20 => "00010110001010010100110001101010",
    21 => "10100011101100110010100111011100",
    22 => "10100001101111010001110011101111",
    23 => "11110011110001100111010110010101",
    24 => "01101111011010011101011111110100",
    25 => "00011111101100110011000000111001",
    26 => "10111000001011101001111100010011",
    27 => "10001101111100011000000010010101",
    28 => "11010110101001010101111100111101",
    29 => "00100010010101111010000111010001",
    30 => "11110010101001100000001001101110",
    31 => "11100110101011111101011101010010",
    32 => "00010100000101100111111111000000",
    33 => "10010000001000101111111001100001",
    34 => "11100110110110111001101111110100",
    35 => "11111001000110111011101011111001",
    36 => "10111011110011011001000101111101",
    37 => "01100011101111011000010001100101",
    38 => "10000110000110111100110001111010",
    39 => "10011010100011100100010011001101",
    40 => "01011001010101010100101010001000",
    41 => "10001000010011111001100011000101",
    42 => "00011000101110010110011100000011",
    43 => "01111010001101010111011010111010",
    44 => "01001110111110001110110011110010",
    45 => "00010101000110100100011010110001",
    46 => "00111010011001111101100011111111",
    47 => "10011101000110101100111000111110",
    48 => "01101011100001000011000011110100",
    49 => "10100100100100001000101111111100",
    50 => "00110111111100111001000001011101",
    51 => "01001111011001001011010101000111",
    52 => "00111010011110110010101111001010",
    53 => "11010001010010111101000001000111",
    54 => "00001010101001100011001110100111",
    55 => "10110110000111001001110010110110",
    56 => "00100110000110111000101000011111",
    57 => "11110101011111110110011111001011",
    58 => "01010100101011010100111011011001",
    59 => "10101110001100111011011101100100",
    60 => "10001100010000011111011100010000",
    61 => "11100101010001010010101100101011",
    62 => "10111111000110000001110000011001",
    63 => "10010101001010000010100011001110",
    64 => "10101111100111011100011000010001",
    65 => "01111100111111000001100111110101",
    66 => "11010111011001001111101111000011",
    67 => "11011011010100100111100001001101",
    68 => "01010010011101110001111111011001",
    69 => "00011000011110000101110110101100",
    70 => "01101110001001001011101011000000",
    71 => "11000110111111111111001000001110",
    72 => "01111101011010001101100011110011",
    73 => "01010011010110010000000100010001",
    74 => "00111111010100110111110010110010",
    75 => "11101110111010101000111001110000",
    76 => "00100110010001001100100000110001",
    77 => "00100110111110001010000101001011",
    78 => "11011000100111101111011110011010",
    79 => "01110101001001011010010111010010",
    80 => "10111110001001111011110111001110",
    81 => "10100001111110111110000011010001",
    82 => "11011110011010101100100100100111",
    83 => "11000110000110000111111010101111",
    84 => "10101011101010000010011001001111",
    85 => "10111001011101011010010110010100",
    86 => "10011101001001001100010000110000",
    87 => "01111101011100010000001110011110",
    88 => "00011100001000101101100010001010",
    89 => "11000110001010100010110101111110",
    90 => "10110000011001001111110011010101",
    91 => "01100011000101110110011010000000",
    92 => "00010010000101101011011000001101",
    93 => "11111101100111100000010111000101",
    94 => "10010001010100010110111110101110",
    95 => "01010011110001101111110101110101",
    96 => "01010101001111111111100110101111",
    97 => "11010100110011000011101001000010",
    98 => "01100011000100111010111110100000",
    99 => "01111001111010010101010011000010",
    100 => "10011010010000010100000110100100",
    101 => "00011100111111101110110011010111",
    102 => "00110001100110111011011000010101",
    103 => "11101000011111000100100111111010",
    104 => "10010100100110000001101010011101",
    105 => "10101100110110101001111110001010",
    106 => "01101111100010110000101111011001",
    107 => "10111011101011101011011000100100",
    108 => "01001011101010000110010000100100",
    109 => "10001000110111100001110111000110",
    110 => "01110101000100100111111110000001",
    111 => "00010000010001110010010001011010",
    112 => "10001110110101101110000111011111",
    113 => "01100101101010101111000110010010",
    114 => "11100101100001111011111100101101",
    115 => "00001110011100111110011010111000",
    116 => "11110110101000100101111101000111",
    117 => "10010111011110110100011000011100",
    118 => "11100100100101001001100011110100",
    119 => "00100000000000111111100011111000",
    120 => "00011000110110001101011011100101",
    121 => "00001101110100111100101101001101",
    122 => "01011100110100001001111010001100",
    123 => "00001010000001011010010010101000",
    124 => "00000010110011110011110101011111",
    125 => "00000101011100101101011010001000",
    126 => "01101111100010001101110110110001",
    127 => "11000010001101000011011000010000",
    128 => "01111010110011010101100101111111",
    129 => "01110000010010100101000100010000",
    130 => "00000111011100110110110111111011",
    131 => "11100000000111100001100110000110",
    132 => "10101010001100010000101101011011",
    133 => "00100110010100111110001010101000",
    134 => "11110111100100001110111110111000",
    135 => "10000111111100100101011111100000",
    136 => "00010011001101100111010000100011",
    137 => "10011000110011011010100101011111",
    138 => "11011111010010001010010010100011",
    139 => "00011000100000000001010101100000",
    140 => "00110101101101110001000001111110",
    141 => "11011001111110011001111011100010",
    142 => "00110011101011001110011011001111",
    143 => "00100011100111111010110111000000",
    144 => "01000100000011001111110010011100",
    145 => "00001110110011110101100100000010",
    146 => "00010010101010000011011010011100",
    147 => "01001001100101100011011111011111",
    148 => "01100110100001101101001000101010",
    149 => "01001011100111101110011001000110",
    150 => "10110110010000011111011000100111",
    151 => "01101110100000011000100001111111",
    152 => "11101001010101110110000101011000",
    153 => "00111001011111110111110011111010",
    154 => "10101010001000100111111111101110",
    155 => "00101010101101111110100000000001",
    156 => "11101111111100100111111001001011",
    157 => "10000101000110010111111010011011",
    158 => "00100000110111110101101111011101",
    159 => "01010010000110011010010101101100",
    160 => "00111100101000110010101100101011",
    161 => "00110000011011001100001100010001",
    162 => "01001111110101100111000011110111",
    163 => "00001100001001001010001110111110",
    164 => "01101001111011010001010101111011",
    165 => "00010100011101010000010100000100",
    166 => "10101011010101001100100000101111",
    167 => "01101001101001110111010111110001",
    168 => "10001010010001011011111101101010",
    169 => "11011101010011000010111110000110",
    170 => "01110101001001101000010101001110",
    171 => "00010100010000011100111111000100",
    172 => "00001100101101011001111001110010",
    173 => "10001000101110000110100010110011",
    174 => "11000010000101000111101010111011",
    175 => "00010010100000010101001011001000",
    176 => "00111011101110110000110010010001",
    177 => "01001110000000110000011110110010",
    178 => "10111100111100010001000011001110",
    179 => "01000001111011101100000010101110",
    180 => "10110001111010110011010101111001",
    181 => "11000111000011010011000111110101",
    182 => "01011001010110100101001100111101",
    183 => "01110001111011000010011100101111",
    184 => "11010011110110111001101011010110",
    185 => "10011000000010000101000111111111",
    186 => "01010111001111000110111001000100",
    187 => "00101110000110110010001110111101",
    188 => "01000101101001010111000000100011",
    189 => "00010001100001110000011100000101",
    190 => "00010001101001011001101010010111",
    191 => "10000110011100011001000011000100",
    192 => "01100110111101100110111110100111",
    193 => "11011000111100100010010010110101",
    194 => "00101110100111000100001111101011",
    195 => "01001010110001011010011011001000",
    196 => "11110001010001001010101100011101",
    197 => "10111101110001110111011100001100",
    198 => "01000010100001111000000010100011",
    199 => "00101110001111110001000100000010",
    200 => "11011111011001010011101110100001",
    201 => "11110010100100011000010011000101",
    202 => "10111010000110100110111111101110",
    203 => "11000100010100111110101111010110",
    204 => "00111111111100001101111111000110",
    205 => "11101111101010011101000011000000",
    206 => "10100011010110100010110110010110",
    207 => "10011010110101110000100100000101",
    208 => "11111010100001111100000011100110",
    209 => "00010111001011010011011110110110",
    210 => "00101001111110101100011001010100",
    211 => "11010111001000000100000001101011",
    212 => "11010011000100001110000100101101",
    213 => "00010111011101011101101110011011",
    214 => "00110000000010101101110010001100",
    215 => "11000111100101110101010100110001",
    216 => "11101100100010100011001111001011",
    217 => "00011100111100000111011110010100",
    218 => "01110010010111111100111011011110",
    219 => "11110010010001100001101010110000",
    220 => "10110111001111011110100111011000",
    221 => "11111000101100110001111100101110",
    222 => "10111000100100000010101111100000",
    223 => "01010110111001000110100110111101",
    224 => "01011100111111010111010100100011",
    225 => "11111000011001010101010001110100",
    226 => "01110110100000111000010001000110",
    227 => "01101110101110100111100011010111",
    228 => "01101001001011010101010111101110",
    229 => "11001010111001000101011110100011",
    230 => "10011100100100100010010100001001",
    231 => "00101000101010000100101010101111",
    232 => "11001100101001001000011011001010",
    233 => "00101111110000001111110010010001",
    234 => "00100110110111010010010110101110",
    235 => "01110001010101010000010001001100",
    236 => "00000011111101110000001010111010",
    237 => "10111000101100110010011011110100",
    238 => "01111101100100100100101110110010",
    239 => "11101111100111110001101101100001",
    240 => "01111101101010010011001000101000",
    241 => "11100001100001111111110001010001",
    242 => "00110111100010100000010010110101",
    243 => "10111101110000010001101111100101",
    244 => "11010110011100101100100110100011",
    245 => "10111001111011111000110100100001",
    246 => "00011011001000010010000001100000",
    247 => "11111100001000010100011110000001",
    248 => "10101000001100001001101000010100",
    249 => "00100110110010011111110011010110",
    250 => "01001101111010010101101101011100",
    251 => "00101101001010001100111101001000",
    252 => "10000010001001110010010010100101",
    253 => "10001110011001111000110010110000",
    254 => "11110101011100111000011011110101",
    255 => "11011010010010010011000100110000",
    256 => "01100110000010110001011111100111",
    257 => "11100111010010010110111110001111",
    258 => "10001100000100111010001010110010",
    259 => "10111110010011000111011100111111",
    260 => "00101101101011111111111100000101",
    261 => "01010101100010110101101100000001",
    262 => "01011010110100111101110000110100",
    263 => "00110000100101101100011010010100",
    264 => "01111101100011101110011010011001",
    265 => "11010010000100100011011000001110",
    266 => "11101111011111111100010010010101",
    267 => "00011101010110001010000000001011",
    268 => "11100101000101101111101110011010",
    269 => "11110001011000000101100110010001",
    270 => "10101001110001101101010011001101",
    271 => "01001101101001110011101110101100",
    272 => "00000111011110101011100001001011",
    273 => "00101101011001110000100101010000",
    274 => "01011001111110110011011010111000",
    275 => "11110110000101001100011101010010",
    276 => "11100011111011111000010011110111",
    277 => "01010000011111000101010100100010",
    278 => "00011101010011001100010011010110",
    279 => "11000001110001111101011101111000",
    280 => "11011000011100111101111100101001",
    281 => "01100110010100111110110101101000",
    282 => "00010011000101010001001011100101",
    283 => "00111001100110101000110011111000",
    284 => "00101111011011001011101000110010",
    285 => "11010010101101101001000100001111",
    286 => "01110110101001000111000101001110",
    287 => "01101001000001010111101110110111",
    288 => "01010101010011100111011111111011",
    289 => "00010001101011011000010010010110",
    290 => "00000010001000000000010110011110",
    291 => "00110110111101001110010001110000",
    292 => "01010011011000100110111000111100",
    293 => "10100100110100101110101111000001",
    294 => "00001000100001000101010101010001",
    295 => "00001011100010101101111010001001",
    296 => "11111010011101001101000011000111",
    297 => "10101000111010111101100000111000",
    298 => "11110101100010110101100101101000",
    299 => "00000101101101011111001000101100",
    300 => "00001101100000010100101110111001",
    301 => "01111110001010111010001010100010",
    302 => "01111000110010100100111111110110",
    303 => "10000010010001001110011010100101",
    304 => "01111101100111011010001101100101",
    305 => "11111101011000100111011010101000",
    306 => "10011011101101001011011100101000",
    307 => "11100101110011010011001110011001",
    308 => "10111011110010001001010010110011",
    309 => "01011111110001100101100001111110",
    310 => "01110001001110101110001010011011",
    311 => "00100101010001010001111001111110",
    312 => "11011101001100000000001011111000",
    313 => "01111001001110011001011100001111",
    314 => "10110000101101110101101111100110",
    315 => "11110111101100110111000000000010",
    316 => "11010111010111000000110001110110",
    317 => "01000010010111100110010010101010",
    318 => "11011101000100000011000011111110",
    319 => "00011110001111110010010001100010",
    320 => "01011000100101011011011010010011",
    321 => "01011010011010110111110101101010",
    322 => "11001111111110001111011000101011",
    323 => "11100011011000011001001100100011",
    324 => "01001010110110001101000001100101",
    325 => "11010000000011100111010011100010",
    326 => "10101110011110010010001010101000",
    327 => "00100111110000110110011001100011",
    328 => "01000011100001001000101000010110",
    329 => "01011110011001001000001000001000",
    330 => "00011111111011001000011010101101",
    331 => "10110010011101001000110110011011",
    332 => "01001011111101110000010010101111",
    333 => "01000111011011101110111110001111",
    334 => "00111001011101100011110110011101",
    335 => "10000011101101010000101000010100",
    336 => "10000001010011111010111100000100",
    337 => "10000110010101100110000111101011",
    338 => "10011110010110010011100010001010",
    339 => "11011101000010100011000000001101",
    340 => "10101100110111111110000010110011",
    341 => "00100101010001011011101111110000",
    342 => "10100010011011000011100001001111",
    343 => "11100111000000100010100100000011",
    344 => "11101110000001100001111111000101",
    345 => "11011010001011001010100001100001",
    346 => "00011011011111101001110100010101",
    347 => "10000101001110110011100110010101",
    348 => "10000001011101000010100001000101",
    349 => "00010000011111001101011101110001",
    350 => "10110010010110000011110100011010",
    351 => "11001100111101100101101000010010",
    352 => "11110010010100100110100100001100",
    353 => "10000100111100001001000101001101",
    354 => "00111101000001001011000100010011",
    355 => "11111001110111011010101010000101",
    356 => "00001111000100110110011001001001",
    357 => "11000101001111011001010100100101",
    358 => "11101100001011001000100011001000",
    359 => "00010111011100000110000011111101",
    360 => "01110001101001100110100100110011",
    361 => "01101000001001010100111011111111",
    362 => "01111110001111100011111101011110",
    363 => "01110100100110101010100000001101",
    364 => "10111010000010101011000110111001",
    365 => "00111010100111001100110110001010",
    366 => "00011001010010010110000100001100",
    367 => "00100000000010101101101011110101",
    368 => "01011010110111111110001110011110",
    369 => "00011100010001110110101110101110",
    370 => "00000110111101100010110110100000",
    371 => "00000001110010010010011001111100",
    372 => "10110101010010000111110010101001",
    373 => "01000111100010010011001010000101",
    374 => "01110011010001100111100111001110",
    375 => "01111011101001111010110111111111",
    376 => "01010000100101101001110011100100",
    377 => "01110010000100011110100101001110",
    378 => "11010001001011011000010110010011",
    379 => "01001110100001110100001111101001",
    380 => "01101011110001000001000011011111",
    381 => "01110111100110110010011000100011",
    382 => "00010000101101110011100100010000",
    383 => "00010000101010010011110000000100",
    384 => "10111100101000010110110101100010",
    385 => "10000011011110111011000101100011",
    386 => "01000011000101011011110111100110",
    387 => "01011001101000010010111011101111",
    388 => "01001100010010111001001110000101",
    389 => "10011001110100110100000000000010",
    390 => "00100100011111101111000001010100",
    391 => "11111001010001111110101100000000",
    392 => "00011111100011110110111000101000",
    393 => "01111101001111010110101100000011",
    394 => "11010101101011011010011111100100",
    395 => "11110111001110101100001110000101",
    396 => "11101110000011101110110111010001",
    397 => "11100100111011101100111100100100",
    398 => "11110011100010010001100101000111",
    399 => "00101011101010001101000110001100",
    400 => "11100101001001111101011110001101",
    401 => "01111100010010011010001010001110",
    402 => "11100111000111001100101000000110",
    403 => "01011111111100110110011111110101",
    404 => "00001000001001110100001101100110",
    405 => "10010110011010101111100000001110",
    406 => "10110000110100011110111011011010",
    407 => "11000011001101110000110101100010",
    408 => "11011010001010000101001110100110",
    409 => "10111110011110000000111100010101",
    410 => "10101001011101011111010001001011",
    411 => "01111101000111101100100110010011",
    412 => "00111101101001001100111100110000",
    413 => "10010110001111010000101111110010",
    414 => "00000011100111011101010101000010",
    415 => "00101000001100101011001100101010",
    416 => "00110000101001000110110011110100",
    417 => "10100111100011101011001101010001",
    418 => "11101101000100011000101111010000",
    419 => "10011000101100010100000100000011",
    420 => "01100111100110010111100000111110",
    421 => "10100001110111110000001011110110",
    422 => "10111110110011110001110000100100",
    423 => "11101000110011001100010000011100",
    424 => "00100101100010101000100011000001",
    425 => "01001000110011010110101101010101",
    426 => "01011100111101111010010111001011",
    427 => "01100110100001010101111100101000",
    428 => "00100111111110011100110110100100",
    429 => "11001011110010100101110101110111",
    430 => "10111110101010000100100010011100",
    431 => "00010100010111010100111110111010",
    432 => "00011000011110010110011001011110",
    433 => "00000111000011011110110010001100",
    434 => "01000011011011100001111001010110",
    435 => "11111010110000111100000101100110",
    436 => "11001110110110110110011010100101",
    437 => "01000011011100101111110110101101",
    438 => "10000001101110001101010010111100",
    439 => "00100110101000011111001010010011",
    440 => "11010011100001001001010011111010",
    441 => "01110110010000111101101010001101",
    442 => "00110101010110111001001011010101",
    443 => "01001011000110001010111111000001",
    444 => "01011001100010111010010011010100",
    445 => "10001000111011010000001101100100",
    446 => "10001010111000000001110111011110",
    447 => "10000111100000001010001100000101",
    448 => "01011001001101100101011000101110",
    449 => "10101000111001000111011001101011",
    450 => "10101110010011011011110100101001",
    451 => "01000111101011000000101100011000",
    452 => "01000000010010101111110000110101",
    453 => "00001010110100111010011010011011",
    454 => "10110111010111101100101010001111",
    455 => "01101001010001110010111001101110",
    456 => "10100000111001001111011100011011",
    457 => "00111011010111111001101001010000",
    458 => "00111100010101000100001010110101",
    459 => "10110011100101011110101001101010",
    460 => "10011101010110110101011101010010",
    461 => "10101110000100111101010011111101",
    462 => "01011001110011010100000011110101",
    463 => "11001011100101001111100101110000",
    464 => "01000100001000110000011110011100",
    465 => "01001111101010000000101110101011",
    466 => "00011000001000011010011110110001",
    467 => "01101111100110011110100010010011",
    468 => "00100010011100110001111110001101",
    469 => "00011010011100000111010011011000",
    470 => "10101011111000110010100001100001",
    471 => "01100100101101010100100110101011",
    472 => "11100011010000101010110001000110",
    473 => "10100011000010001010100101101101",
    474 => "10100110100011010010111000010000",
    475 => "00110101011101101101011010001000",
    476 => "00010011001000011000000110101010",
    477 => "01101100001000111111101010010110",
    478 => "10011001000111110010001110001101",
    479 => "00011111111100100101100111000110",
    480 => "10101100001100100110001111100011",
    481 => "11001111101100101110111111101111",
    482 => "10000110111011100111110000110101",
    483 => "00011100110000001010111101111111",
    484 => "00111001101110100110011110110101",
    485 => "00000011001100111000010111100011",
    486 => "10111010111010001100011110100111",
    487 => "10110010011001011010111110010010",
    488 => "00000111111111011011001110001001",
    489 => "10111101110000100110001011101101",
    490 => "00101100000011001110110011011100",
    491 => "11110010011100110110011100000000",
    492 => "11010110110000111110010011111011",
    493 => "00101100000111010011000100101010",
    494 => "00010110010100000101010110011110",
    495 => "01001101001001010011001110110110",
    496 => "00111011101010011111000001100010",
    497 => "10000110110101101100010100011101",
    498 => "01011100001001001111110000101111",
    499 => "11101011111110100000100001011101",
    500 => "11011010110010001001100011111001",
    501 => "01111011011111001111001111111110",
    502 => "01010111000101100101110111001111",
    503 => "00110011110111001101010010010001",
    504 => "10000011010100001111110010010101",
    505 => "10001101100111101111001011110111",
    506 => "11100100110110000111000011110100",
    507 => "11101110100011000101011111110111",
    508 => "11011110101010011011101110010010",
    509 => "10101011011111110101111001111100",
    510 => "01100110101110010001010000010010",
    511 => "10110111011111001100101010111001",
    512 => "10010101011111001011010111011111",
    513 => "11100100111110110111000100001111",
    514 => "11100001111010110000010001110100",
    515 => "10000111100000010001010111110011",
    516 => "01000000001000110000011110101101",
    517 => "01010010011001001111111000010001",
    518 => "10110000111000001010110110000110",
    519 => "11110110010011010111011011010110",
    520 => "01110111111000010000101000100001",
    521 => "11100011100011111001001110001100",
    522 => "10000011111111101100001111001100",
    523 => "10011000010101011101000100001000",
    524 => "01101100110001010111010010101001",
    525 => "01010111101000101001000010010011",
    526 => "00111100011110011100000110111010",
    527 => "11110101111000011000110100110011",
    528 => "11001101011100101110101100100100",
    529 => "01000011100110000010100110101000",
    530 => "00101011110100100111011110101111",
    531 => "01101100000100011000110100001101",
    532 => "01001110000101110100100110010000",
    533 => "00000011001011101110010011011001",
    534 => "01000100101110000101110111000100",
    535 => "00110011001010011010000100110010",
    536 => "11111101011010001100010110000000",
    537 => "00011001010100101110001011111110",
    538 => "01101000110101010010000001000111",
    539 => "01100100000100000000100010110000",
    540 => "11110101011111011110001110001011",
    541 => "00101001000110010001110110101100",
    542 => "01001010110100011111010010010100",
    543 => "10000011111011100001110011100011",
    544 => "11111001110101111010100100100010",
    545 => "01000111101000101100111101010100",
    546 => "00010010100111111000011000101110",
    547 => "10010001100111111010000000101101",
    548 => "01110010001010101110011110000011",
    549 => "11011111101011101100011011011010",
    550 => "00001110010010101110000010111010",
    551 => "01110011011111001010110100101101",
    552 => "10101001100100011001110011001111",
    553 => "00001101000110110010111110001100",
    554 => "00111110011110000100010000110011",
    555 => "11101000000000010101001000000111",
    556 => "10101100110111011101000101111111",
    557 => "11100101111011011100110100001100",
    558 => "10110000000101010001101010010110",
    559 => "10001111111101001010010111010000",
    560 => "10110001011000100011000001111111",
    561 => "01001111100101101110010010001101",
    562 => "10001011010010111101000110001010",
    563 => "00100100101110001000011001110001",
    564 => "11110110000001010000100111000110",
    565 => "10110100010110011111111001010110",
    566 => "10010111001111111011010101010111",
    567 => "10010000000000111001000010111011",
    568 => "10110100101001100011101110110011",
    569 => "01010011001110000000111100111101",
    570 => "10001110010010011111100010000011",
    571 => "10100111000101001010011110101001",
    572 => "11001100010100111101000011111011",
    573 => "10110010110101111001000000011011",
    574 => "11110110110111100101111010101001",
    575 => "10100110010101011010111101001010",
    576 => "00011010011000111010101100010100",
    577 => "11101100010000100100010111011011",
    578 => "11010111001000110001100010010111",
    579 => "10100011001001100011010110101101",
    580 => "10010101011000100001100110010111",
    581 => "01010001011110000000110011011101",
    582 => "01101101011100110010000100011001",
    583 => "10100111000110111001101100100100",
    584 => "11111011111001001001000110011111",
    585 => "01001000000011000010000001101111",
    586 => "11011011001100101011011110000111",
    587 => "11000100101000010100111000101101",
    588 => "10111101101011111110011001111001",
    589 => "01111010010100011010010101011001",
    590 => "01100000111000111001000101010011",
    591 => "11111101110000110000111000101101",
    592 => "11110111100011101011011110000000",
    593 => "10000101001011101100110001000111",
    594 => "01111000011010010111011111011101",
    595 => "00111001100100101010000000001010",
    596 => "10111000001000100111011010111110",
    597 => "00101011101111010111001010100001",
    598 => "11100111101100001111000101111010",
    599 => "01000011101000010010101100001110",
    600 => "00100001000010010101000010010111",
    601 => "10101011110011011110010110110101",
    602 => "00000110100100001111110000001011",
    603 => "01001110010011010001111001001111",
    604 => "01011011011001100011000101011101",
    605 => "00011100010101000111010000010111",
    606 => "00101111001100101010111011100001",
    607 => "11110100010100000110110010011011",
    608 => "00111011000000001100011000100010",
    609 => "10110011101100100011011101111101",
    610 => "01010000001001100001001000001000",
    611 => "10101011001010101001010101101010",
    612 => "00010100010010101001100010101010",
    613 => "00111111000001010101110101101100",
    614 => "10101001110000010001010111010110",
    615 => "11011111100100010000110101000011",
    616 => "00001110010100111101001111111000",
    617 => "01000111000001100110111010001100",
    618 => "11111011110011100010011011011110",
    619 => "11011001001001011011001010010001",
    620 => "01011101111100100101000010000011",
    621 => "10010011011111100001101011101100",
    622 => "00001111100100011010100011110000",
    623 => "00110011111001100110010111001010",
    624 => "10000001010011011100000001101011",
    625 => "01111101111111001010110100011001",
    626 => "01010100110111010111010011001110",
    627 => "01011001101111000101101100111001",
    628 => "11100101001000111001011110011101",
    629 => "00011011011010000100000100100000",
    630 => "11110100100110101100011011010011",
    631 => "11010000000100111001011111011100",
    632 => "00111110101000001110010100100101",
    633 => "01010000111101001100001000111010",
    634 => "00100011000101100001011011110110",
    635 => "00001101010000001011111001011110",
    636 => "10111100000011000001001000100110",
    637 => "10111110011000101011100101101010",
    638 => "11100111011001001101011001101000",
    639 => "01010111100010110001010100110111",
    640 => "10010001001001000100110001001000",
    641 => "10001110100010001100011000000100",
    642 => "00010101100100001001011101111101",
    643 => "10000011101000100110000000101011",
    644 => "00111000011010000111000011111101",
    645 => "10111111011010001101001111111111",
    646 => "11001000110001101011011001101000",
    647 => "01101000101001000110110100110011",
    648 => "11011011010111100010101010010110",
    649 => "00011111001011100011001101000011",
    650 => "11101000100000000100001000101111",
    651 => "00110101000010000111001101101111",
    652 => "01001001010000010101100011110111",
    653 => "00010100011111101100110001001001",
    654 => "10110011000110111010011010101111",
    655 => "00010110000001111011001011100000",
    656 => "10011000011100100110101110001001",
    657 => "00101111001000001001101001111101",
    658 => "00110011001010001000100101111001",
    659 => "10101000101101110011001000101001",
    660 => "01010001110011011001101111110011",
    661 => "10011000100101000011001001001011",
    662 => "01110111100111000111001000001001",
    663 => "00100001111110111110110111101101",
    664 => "00111010110100011100111011101100",
    665 => "11010001011011101101111000110000",
    666 => "11101101100110010001001011011010",
    667 => "11000111110111100110010101111000",
    668 => "11111001111000100111111001111100",
    669 => "11100111100000001001101100110001",
    670 => "11001000011001110001001101000101",
    671 => "11110001001111100001100000100111",
    672 => "00100010000110001100011011110111",
    673 => "00001110110111001000000111011100",
    674 => "01010011001000011010110101001100",
    675 => "01000000110100100100101011101010",
    676 => "00011111101100111011101000101111",
    677 => "10111111100000111001101110011111",
    678 => "01011010100111110001110010110100",
    679 => "01101010010010101100100011011011",
    680 => "10100010101010011010101011000110",
    681 => "10111000110000101111110010111111",
    682 => "01000010001100001111100010101010",
    683 => "11000111000111010010100101110010",
    684 => "01011100111111101001001111111100",
    685 => "01101001000100011001110001010110",
    686 => "00101100001001100001001010110110",
    687 => "00000110001111110010011000010011",
    688 => "01111010101011100110011100100001",
    689 => "00100011100000000010101000011101",
    690 => "11001100101011110101101111110101",
    691 => "11110010101111110101110110101101",
    692 => "00111101101110001111001000111101",
    693 => "00000011101100110100001001100000",
    694 => "10010011110000101000001011100001",
    695 => "00101101110010001111101010010101",
    696 => "00101001101101111011001001000111",
    697 => "01000110101011101110101101001000",
    698 => "01100111001011010101100110001111",
    699 => "10100111111111000010001000011101",
    700 => "10111100011010011101100101011110",
    701 => "11101001100100011001010011001100",
    702 => "01101011010111010111001011110001",
    703 => "00110110110011101100010111000001",
    704 => "10000100111011000110001011010010",
    705 => "00110011110110111110111010000000",
    706 => "00111110101000010110010011101010",
    707 => "10111101111111101101010011110100",
    708 => "01011000110111100100010110000001",
    709 => "00010100101100100110011000011100",
    710 => "00101111101100000010001010010101",
    711 => "00100011000011001111011000001010",
    712 => "10101001000001110101100000000101",
    713 => "01000101010100000111111111010010",
    714 => "11110111100001111111011000001101",
    715 => "11010100011000001001111100011111",
    716 => "01111110010110100110000001100111",
    717 => "10011100100000011011101110000000",
    718 => "00101101110000101110111011010010",
    719 => "01001111110000111010110101101110",
    720 => "10101101100111110111000100100000",
    721 => "00000100010010110001000001110000",
    722 => "00101010001110101110100000100011",
    723 => "01101000100110110010110100110101",
    724 => "00000011111110111111110010111110",
    725 => "11101111101110011111011000001000",
    726 => "10111111110010001111010000000010",
    727 => "00001101000100111111010000101111",
    728 => "11111100100000101100110101100101",
    729 => "11111001000001001111110110011111",
    730 => "00111111101100010001010111111001",
    731 => "10100111111111001001001011011101",
    732 => "10001011010101111101000010101101",
    733 => "00100111110000110100100110111100",
    734 => "10010111110011101100111110011111",
    735 => "11101011110010100001000100100111",
    736 => "11111011001001101001001100100001",
    737 => "00110001101011110001011011001101",
    738 => "00110010010111110000011100000001",
    739 => "00101000011110101010100011101010",
    740 => "10010111100101111101011101010011",
    741 => "11101010000001110010001100010010",
    742 => "10101010111110111000101100000100",
    743 => "01000000001100010001011101011100",
    744 => "11001001011111111000101101000111",
    745 => "00011011100010010001101111011011",
    746 => "00000110100110111011000110111101",
    747 => "11000111001111000001011110100101",
    748 => "00001000000000111111110100010110",
    749 => "01001011000011100100000111101101",
    750 => "01100110100001100101100010010001",
    751 => "11100101010000010000110101110100",
    752 => "10100110111011010111010010101100",
    753 => "10000111000011100110011011110111",
    754 => "00110001001110100110100001000011",
    755 => "00001111101001110111111101101100",
    756 => "01000111101111011010111011010011",
    757 => "10100000001100110000101011101011",
    758 => "11110000110010011011100111000100",
    759 => "10011010001101111001001001000001",
    760 => "10011001100110100011011101000110",
    761 => "11000011011110011110011001010000",
    762 => "11111001010001100101110011010110",
    763 => "00110010001010010110101101110001",
    764 => "01111001101101010101111101011000",
    765 => "00100001000111010010011010100010",
    766 => "00110100000100000000000001110011",
    767 => "11000001111010001010001110011111",
    768 => "10011101010011100101100001011100",
    769 => "10110100010010011111000011010001",
    770 => "01111000100000000001101001111100",
    771 => "00010111010110110000000000111010",
    772 => "00111101101000000001001011000000",
    773 => "10110010111101110000001100101100",
    774 => "00010111111100100010110101110101",
    775 => "11101000101100110001000110001111",
    776 => "10000010111011110100001110001110",
    777 => "01010001110000100100110111000011",
    778 => "10110110111000101111010111010110",
    779 => "11111101011111111111101001010101",
    780 => "00000001001000110110011010010011",
    781 => "10010000110101000000110100011111",
    782 => "00100100111110110101010100010101",
    783 => "00010000001100001101110000100101",
    784 => "00011011101100111011101101011001",
    785 => "10010000110100100110111000010101",
    786 => "00001000011011000011110100111000",
    787 => "01010100011100011001111100101110",
    788 => "01011111101110110111100101111100",
    789 => "11110100011101100001110001111100",
    790 => "01010100100101110011011111001011",
    791 => "00101001001110100000101110101101",
    792 => "00001001010101100010010111101111",
    793 => "11010011101111000001101111000110",
    794 => "11110000110100010111000011110111",
    795 => "11101111110110010011011100010110",
    796 => "00110101001111101110000000111101",
    797 => "01010100011000100010111011011001",
    798 => "01010111000111100011100110100001",
    799 => "10001001111010101000100101011101",
    800 => "10000100010010011100000000001100",
    801 => "10010000000111100001011000001001",
    802 => "11011000011000110001011010001101",
    803 => "01100000001001000000000110011000",
    804 => "11100111100001110011011001110111",
    805 => "10101010000000100110000100011001",
    806 => "00001100010000011011010011000010",
    807 => "00001011101111011001101110011000",
    808 => "01110011100100011010001011001110",
    809 => "00110001001110011110011010101000",
    810 => "10001010101100010010011101111000",
    811 => "11100110000010001001000111100000",
    812 => "10110101111001111010100111101110",
    813 => "00000101010111111100010000100001",
    814 => "00101010100000001010101011101111",
    815 => "11110100111101101000101101000110",
    816 => "00100001101000010001010000011000",
    817 => "00000111100001011100101000111010",
    818 => "11110100111011100011000011011010",
    819 => "11000110110111010101110110110011",
    820 => "00011100011001010000010100110111",
    821 => "01101101001101101010100101111110",
    822 => "10100100001110000100010111010100",
    823 => "10001000101001001000101010000101",
    824 => "00000011100110011111001101010111",
    825 => "01111100001011001111110001101100",
    826 => "11011010111100011000111011110000",
    827 => "11001110001110110010001010001110",
    828 => "10011100101000000100111100001001",
    829 => "10011101110111110001110001101110",
    830 => "01100010111001010011010000101101",
    831 => "11110101111010110110010011111000",
    832 => "00010111111010100100100100001001",
    833 => "11100101000110101111101100000110",
    834 => "11101001010011011110000100111100",
    835 => "00110110010001111000111101101110",
    836 => "00101010001001101011101000111010",
    837 => "11001111011110001100111111010001",
    838 => "11110010010010011011110111100101",
    839 => "01101100101010011011010111110001",
    840 => "01100001010111011101111000000000",
    841 => "11010000101011000100100010100101",
    842 => "01011000011101000111110110111111",
    843 => "10000011001100111110011100111101",
    844 => "00110100011011011001000110101010",
    845 => "00001001001010010100000111100111",
    846 => "11101010100111110110001110110100",
    847 => "10100111110010100010010111010110",
    848 => "10101101111011000000010011010111",
    849 => "00101110100100011010011101000101",
    850 => "00001110011001010010000100011001",
    851 => "01101101101111100111000011001110",
    852 => "00111111010110010000101111110110",
    853 => "11101011010101110010000000011010",
    854 => "10010000010010100000001111001111",
    855 => "00100000000110011000010000110000",
    856 => "10011111100111000001101011110000",
    857 => "10100001010000001110001001011110",
    858 => "01011110000100100110010010000111",
    859 => "11101110011001000011001011100010",
    860 => "10001010100011011110010100000111",
    861 => "00111100110110001110110011010100",
    862 => "10011000101000001111111110111001",
    863 => "11011110010101110001111101011111",
    864 => "01110001100010000011001110000110",
    865 => "11011101110001101110101010100111",
    866 => "11110001110000011111110101011000",
    867 => "00111000011110010010111111110110",
    868 => "00001000101111001001110000011100",
    869 => "11100010101111011101001100101101",
    870 => "01111011110100010010011000100000",
    871 => "10001010101011101000000110111100",
    872 => "01110011100111010010010000110110",
    873 => "00010011011111011101100111000001",
    874 => "01010000011001000010110110110110",
    875 => "11100100001011110111111011101110",
    876 => "11111001011011111000000101101100",
    877 => "01010000000111110101101101111101",
    878 => "10000101101010110111111001101101",
    879 => "01011000100111011000010110111101",
    880 => "10111011010111110100000110000100",
    881 => "01110111001000010000011010010011",
    882 => "10000001111010011100101111011110",
    883 => "01011110001111000100100000101110",
    884 => "01010011011010101000011010011111",
    885 => "10100011101011010000011111100110",
    886 => "11000011110100010111001010111000",
    887 => "11101010101010001110110111010000",
    888 => "01011010010010101110110110111101",
    889 => "00001001000111100001111110101011",
    890 => "10000101101000010010111000110101",
    891 => "00001110010101100000101001011101",
    892 => "10001011100010001101011011010001",
    893 => "00000100001101110000010010001110",
    894 => "00001011001101010011101010111110",
    895 => "00011010100010101100110011110011",
    896 => "01101100101101111000010011110011",
    897 => "00110001111100000111011111100100",
    898 => "00100111000110110000000011001111",
    899 => "10001011111011011110100001111101",
    900 => "01010100100101101010101101000110",
    901 => "01111001001000111001001001011100",
    902 => "10000111001011011111001000101000",
    903 => "00111101011001100110000010101100",
    904 => "11111110000111011001101110010001",
    905 => "11111101100110011011000001110001",
    906 => "10110110111001111000101010010001",
    907 => "11011001011111110101001101111000",
    908 => "00011111111100010100001110011101",
    909 => "10100110100101101011110111110001",
    910 => "10011101010011001001111000011100",
    911 => "10101101011111001011111110110001",
    912 => "11011101100101100010001110111001",
    913 => "01010100111101111111000000110001",
    914 => "01100100110010000011011000011100",
    915 => "01001111011110010010110101000111",
    916 => "00110000101001010011001111100111",
    917 => "11111000100111100111101001111010",
    918 => "00011100000010110011111111000001",
    919 => "11001000000111110011011111100011",
    920 => "11110011011101000001000000010011",
    921 => "00011101111001111010010100011100",
    922 => "01010001101010001010001100100111",
    923 => "01101100110010111111110000001000",
    924 => "11010101000111010101000010100010",
    925 => "00011100110000000110010100011111",
    926 => "01010100100001000100010011011110",
    927 => "11111100011011100001000111010010",
    928 => "00101001101010100101110001101010",
    929 => "10110110110010111000110100101000",
    930 => "00110010010010111101101010110101",
    931 => "01000111110100010111001111101010",
    932 => "11001110111000010111101000010011",
    933 => "00011010110001000011010010101100",
    934 => "01110110011101001100100110010010",
    935 => "10000101000101011001010100101110",
    936 => "00101000100111000101010011100111",
    937 => "00010100010001000111010001001011",
    938 => "00011010011001000011001011100010",
    939 => "11101011110111101101111011010010",
    940 => "00010100011100110010101001001100",
    941 => "11100001111010110111001001000110",
    942 => "01010010110111000110100011000111",
    943 => "00011011000100011101011111000110",
    944 => "00101111101111111000011000011011",
    945 => "10001010111110010101011110111100",
    946 => "11011000001000100001111101011110",
    947 => "11000100111111000110111101101101",
    948 => "00010011001110101011101000010010",
    949 => "00010001111100000101001101001101",
    950 => "01000010101001000001000010101100",
    951 => "11110011100110000101110101001011",
    952 => "10111010000000110010001011000101",
    953 => "11100101100001010101110110100010",
    954 => "10001000111011010100000111101001",
    955 => "01000011111010001101100100101111",
    956 => "01011010000000111000000001100110",
    957 => "10000110010101111101101101100000",
    958 => "00000100001011011100111110001110",
    959 => "00101001011001101010111001100111",
    960 => "01110011010001110001100000011000",
    961 => "10010101111110001011011001111110",
    962 => "00000111001010101101000111001110",
    963 => "01110010011011001101000011101111",
    964 => "10111010101101011100101000001000",
    965 => "00100100000101010000111110000101",
    966 => "00011011011000110000110010110111",
    967 => "11101000100110100100000001000111",
    968 => "10011111100010100011111001100110",
    969 => "10101001110011011000010100100111",
    970 => "00011111100000111101101001011110",
    971 => "11000101110101111110110010000101",
    972 => "00010011100010101010100111010000",
    973 => "10100110011001110100001111111010",
    974 => "01101101100110010111101100010011",
    975 => "01001011101001011100111100001111",
    976 => "00000100001011011111100010000100",
    977 => "10101100010010011100101010100110",
    978 => "00111100100100111010101101111100",
    979 => "10100101101111100101011000110111",
    980 => "00100011000100111011111111010010",
    981 => "01110100101000110101000000111100",
    982 => "11100001100000001101001010010001",
    983 => "00010011110111001111110000001010",
    984 => "10101011010111010010111001110001",
    985 => "00101001100000101001000101001011",
    986 => "10101011011000001101111110001100",
    987 => "11000100011010000110001110011100",
    988 => "10111011100010100100010110111101",
    989 => "01010110101001000000001011000010",
    990 => "10111010100111011001100111110111",
    991 => "00001010000001000101001111111011",
    992 => "00000011111010000101011101011111",
    993 => "01001010001001000101110011010010",
    994 => "11010101000001001011101000111011",
    995 => "10110111110001010111100001101000",
    996 => "10111001101101100001100011001101",
    997 => "10110110100011110100011010011010",
    998 => "10001001101001100101100100101100",
    999 => "10011100010000011111110001011010");

  constant ans_lut : lut := (
    0 => "00001101000100110111011011011110",
    1 => "10000100001100010111101101001010",
    2 => "10110011000111001001011010011110",
    3 => "00010000110110001001001010110000",
    4 => "10011101111001110000100111100010",
    5 => "01001000011101100101000010101110",
    6 => "00101110011001001010011001010000",
    7 => "00111001010101010010001100100000",
    8 => "11100011101001010001100101110010",
    9 => "11110000111010111111110010010000",
    10 => "11011011100100100011011010100010",
    11 => "11000000001001101000101001100100",
    12 => "11001110011110100100010101111010",
    13 => "01010100001001010011100101110100",
    14 => "10101111110110100100001110111010",
    15 => "00000011011110011110100010111010",
    16 => "00010110000110010011100010010100",
    17 => "01110101111011010000110010011010",
    18 => "00111101000000100010111110101010",
    19 => "00000100010111110100001001110010",
    20 => "01101000110000011000110100110110",
    21 => "11011011001101101110010011110100",
    22 => "11011101001011010100010110100110",
    23 => "10001011001001010001110010101000",
    24 => "00001111100011000010000010111110",
    25 => "01011111001101101101111001110100",
    26 => "11000110101110111010011011010110",
    27 => "11110001000001111010111100011110",
    28 => "10101000010001100010010110101110",
    29 => "01011100100101111111011001101010",
    30 => "10001100010001010110001011100110",
    31 => "10011000001110100101100110100000",
    32 => "01101010110110011011101010011110",
    33 => "11101110110010010000100111011010",
    34 => "10011000000101010011010111100100",
    35 => "10000101110100100110101000111100",
    36 => "11000011000111110110011011101010",
    37 => "00011011001011001110011100001100",
    38 => "11111000110100100101001010011000",
    39 => "11100100011001100101001100011000",
    40 => "00100101100110011010000101100000",
    41 => "11110110100111011101100000110000",
    42 => "01100110001100001011110101101010",
    43 => "00000100101101001001001101110100",
    44 => "00110000000000111010001101000010",
    45 => "01101001110101000110010111111010",
    46 => "01000100100011010101010110001110",
    47 => "11100001110100111010110000000000",
    48 => "00010011011101111110001000100000",
    49 => "11011010011000101011000111011100",
    50 => "01000111000001101000100100010110",
    51 => "00101111100011110100011000111010",
    52 => "01000100100000100111010111111110",
    53 => "10101101101000001100011000111100",
    54 => "01110100010001010010100001101110",
    55 => "11001000110100010011101011110010",
    56 => "01011000110100101010110001010010",
    57 => "10001001100000000100110001001000",
    58 => "00101010001111010001001011100100",
    59 => "11010000101101100101010011101110",
    60 => "11110010101010001111000000001000",
    61 => "10011001101001100011000101011100",
    62 => "10111111110101110110110001100010",
    63 => "11101001110000101101110011011010",
    64 => "11001111010011111011000010011100",
    65 => "00000010000000011111101010111110",
    66 => "10100111100011110001101000100010",
    67 => "10100011100110111011000010010000",
    68 => "00101100100001001001100011011110",
    69 => "01100110100000111110111100110100",
    70 => "00010000110001101110101110000110",
    71 => "10111000000000000000011011111000",
    72 => "00000001100011001011101000110010",
    73 => "00101011100101110000000001110000",
    74 => "00111111100110101111000011011110",
    75 => "10010000000010111011001110110110",
    76 => "01011000101001101000010011110000",
    77 => "01011000000000111100101101010000",
    78 => "10100110010011100010000101101100",
    79 => "00001001110001011101000101000000",
    80 => "11000000110000110101100100101000",
    81 => "11011101000000100001100000111010",
    82 => "10100000100010111001000011001000",
    83 => "10111000110101101110000100011110",
    84 => "11010011010000101101111111000000",
    85 => "11000101100001010110010100010010",
    86 => "11100001110001101110000000100100",
    87 => "00000001100001111111010101110100",
    88 => "01100010110010010011100010010000",
    89 => "10111000110000001000110100111010",
    90 => "11001110100011110001100101110110",
    91 => "00011011110110000110111011000110",
    92 => "01101100110110010110110000101100",
    93 => "10000001010011110101110011100010",
    94 => "11101101100111000111010101001000",
    95 => "00101011001001001010101111101000",
    96 => "00101001101010101011000001001000",
    97 => "10101010001000000111001011001100",
    98 => "00011011110111011110000001001000",
    99 => "00000101000011000110111110000100",
    100 => "11100100101010011000111010011110",
    101 => "01100010000000001000101000101000",
    102 => "01001101010100100111000011011000",
    103 => "10010110100000011110000111111110",
    104 => "11101010010101110110111001111100",
    105 => "11010010000101011110001000101010",
    106 => "00001111011010111010100110011100",
    107 => "11000011001110111000111000001110",
    108 => "00110011010000101001100000110000",
    109 => "11110110000100111000011010111110",
    110 => "00001001110111111010110011011110",
    111 => "01101110101001001000101111000010",
    112 => "11110000000110000111111000100110",
    113 => "00011001001111111011000001011100",
    114 => "10011001011100010110001111111110",
    115 => "01110000100001100101100101111000",
    116 => "10001000010010011100111011010110",
    117 => "11100111100000100110100001010100",
    118 => "10011010010111001000001111100000",
    119 => "01011110111110000100101101001000",
    120 => "01100110000101110001110111001110",
    121 => "01110001000110101011011101011110",
    122 => "00100010000111010001001000011110",
    123 => "01110100111101010011000010110000",
    124 => "01111100000111100001110111001100",
    125 => "01111001100001101111000000001110",
    126 => "00001111011011110110101010101010",
    127 => "10111100101101011101010011000100",
    128 => "00000100000111111001001001100000",
    129 => "00001110101000011111011011000100",
    130 => "01110111100001101001110000011000",
    131 => "10011110110011110100001011111010",
    132 => "11010100101110010001010101100010",
    133 => "01011000100110101010011001001110",
    134 => "10000111011000100001010111011010",
    135 => "11110111000001110011011010010100",
    136 => "01101011101100111001100010101000",
    137 => "11100110000111110101010001100110",
    138 => "10011111101000110101000010011010",
    139 => "01100110011111111101010101000110",
    140 => "01001001001100101111111101000010",
    141 => "10100101000000110100010101101100",
    142 => "01001011001111011000010010101010",
    143 => "01011011010011010011011001001100",
    144 => "00111010111010000110101101000000",
    145 => "01110000000111100000100010111010",
    146 => "01101100010000101100110011100000",
    147 => "00110101010110100010001011001110",
    148 => "00011000011100110000110001011100",
    149 => "00110011010011100011011111100110",
    150 => "11001000101010001111000011010100",
    151 => "00010000011111001111100001001100",
    152 => "10010101100110000010001111100100",
    153 => "01000101100000000100000110100110",
    154 => "11010100110010011010011001001010",
    155 => "01010100001100100010110101111110",
    156 => "10001111000001110010000100100110",
    157 => "11111001110101010111101011011000",
    158 => "01011110000100101011010010100010",
    159 => "00101100110101010100010011101000",
    160 => "01000010010010001101001010101010",
    161 => "01001110100010100110011010001100",
    162 => "00101111000110001100111001110010",
    163 => "01110010110001110000011101010110",
    164 => "00010101000010100011011001110010",
    165 => "01101010100001011011110001111010",
    166 => "11010011100110011111111101111110",
    167 => "00010101010000111010110100000000",
    168 => "11110100101001011011010011000100",
    169 => "10100001101000000111101100111010",
    170 => "00001001110001001100011111000100",
    171 => "01101010101010010001001001001000",
    172 => "01110010001101000110101111111000",
    173 => "11110110001100011011000100100110",
    174 => "10111100110111001011000011000100",
    175 => "01101100011111010110000101011100",
    176 => "01000011001011110010111100011000",
    177 => "00110000111110100001010001111100",
    178 => "11000010000001111110111000000100",
    179 => "00111101000010010011111100100010",
    180 => "11001101000010110101000010000010",
    181 => "10110111111010000001001101110010",
    182 => "00100101100101100001011010001100",
    183 => "00001101000010101100000111101010",
    184 => "10101011000101010011011010100110",
    185 => "11100110111100000110000000000010",
    186 => "00100111101011011110011001000010",
    187 => "01010000110100110011011101010110",
    188 => "00111001010001100001000101110000",
    189 => "01101101011100101010110100111000",
    190 => "01101101010001011101111010101010",
    191 => "11111000100001111010011000001000",
    192 => "00011000000001001111011110101100",
    193 => "10100110000001110101001100100100",
    194 => "01010000010100011011000111010100",
    195 => "00110100001001011100100101101010",
    196 => "10001101101001101001110110010000",
    197 => "11000001001001000100011110001010",
    198 => "00111100011100011101001101100110",
    199 => "01010000101010111000000000100100",
    200 => "10011111100011101111001001000000",
    201 => "10001100011000010010111001000110",
    202 => "11000100110101000010110101000110",
    203 => "10111010100110101001111110011100",
    204 => "00111111000010000000100110110010",
    205 => "10001111010000001111011001100010",
    206 => "11011011100101100011000001110010",
    207 => "11100100000110000110001001100010",
    208 => "10000100011100010110000011110000",
    209 => "01100111101111010010110000100100",
    210 => "01010101000000101010101011000010",
    211 => "10100111110011000111101001110110",
    212 => "10101011111000100010110010001100",
    213 => "01100111100001010100011111000000",
    214 => "01001110111010111111100111100000",
    215 => "10110111010110001000011110000110",
    216 => "10010010011011010001101000000100",
    217 => "01100010000010000100010010100010",
    218 => "00001100100100100110100101000000",
    219 => "10001100101001010110100001100110",
    220 => "11000111101011001000101010110010",
    221 => "10000110001101101110111111100000",
    222 => "11000110011000110100100011111000",
    223 => "00101000000011110111010110011100",
    224 => "00100010000000010100100010110010",
    225 => "10000110100011101110001011001000",
    226 => "00001000011110010010011110011000",
    227 => "00010000001011111011100111011110",
    228 => "00010101101111010000101100101010",
    229 => "10110100000011111000000011111100",
    230 => "11100010011000000011011101010110",
    231 => "01010110010000101011010110100100",
    232 => "10110010010001110010101001011100",
    233 => "01001111001010011100101101001110",
    234 => "01011000000101000010110000111100",
    235 => "00001101100110011101010000001010",
    236 => "01111011000001001010100010000010",
    237 => "11000110001101101110011111101010",
    238 => "00000001010111111111110000010110",
    239 => "10001111010011011111001100010100",
    240 => "00000001010000011010101101000000",
    241 => "10011101011100001111011101110100",
    242 => "01000111011011010110101011101000",
    243 => "11000001001010011010111111000010",
    244 => "10101000100001101111011100111010",
    245 => "11000101000010001100101000000100",
    246 => "01100011110010110101111001000000",
    247 => "10000010110010110010110011101110",
    248 => "11010110101110011000110000011010",
    249 => "01011000001000100011101001001100",
    250 => "00110001000011000110101110001100",
    251 => "01010001110000100001110010110000",
    252 => "11111100110001000000110000101100",
    253 => "11110000100011011000010000100010",
    254 => "10001001100001101000111001001100",
    255 => "10100100101000101101111010000010",
    256 => "00011000111010111001010100110010",
    257 => "10010111101000101010110000010110",
    258 => "11110010110111011111001110110110",
    259 => "11000000101000000100001011110010",
    260 => "01010001001110100010111110010110",
    261 => "00101001011010110010001111000000",
    262 => "00100100000110101010101100001000",
    263 => "01001110010110010101010001010110",
    264 => "00000001011001010100111001010110",
    265 => "10101100111000000001110101000000",
    266 => "10001111100000000001110110111110",
    267 => "01100001100101110100010000010010",
    268 => "10011001110110010000100000000100",
    269 => "10001101100100100000111010111110",
    270 => "11010101001001001100110110010100",
    271 => "00110001010000111111000100101110",
    272 => "01110111100000101011001000010110",
    273 => "01010001100011011101010010011010",
    274 => "00100101000000100111000001010000",
    275 => "10001000110111000011111100101000",
    276 => "10011011000010001100111010101110",
    277 => "00101110100000011101110001000000",
    278 => "01100001101000000000011000111010",
    279 => "10111101001000111111100001000100",
    280 => "10100110100001100101110110100000",
    281 => "00011000100110101001111001111000",
    282 => "01101011110110111100111110000100",
    283 => "01000101010101000000010101100100",
    284 => "01001111100010100110101110111100",
    285 => "10101100001100110111110000110010",
    286 => "00001000010001110100010001100000",
    287 => "00010101111101010111101111100100",
    288 => "00101001100111101011010011110100",
    289 => "01101101001111001101100001010100",
    290 => "01111100110011001100010110011100",
    291 => "01001000000001011100111001000010",
    292 => "00101011100100001011011100100010",
    293 => "11011010000110110101101101011000",
    294 => "01110110011101111001111000000100",
    295 => "01110011011010111111011010000000",
    296 => "10000100100001011101100100000010",
    297 => "11010110000010101111000001011100",
    298 => "10001001011010110010011001110010",
    299 => "01111001001101000001100011110000",
    300 => "01110001011111010110111100110100",
    301 => "00000000101111101110101010011110",
    302 => "00000110001000011111011110101000",
    303 => "11111100101001100110101100110010",
    304 => "00000001010011111101111001001100",
    305 => "10000001100100001011000111000100",
    306 => "11100011001101010101001011100000",
    307 => "10011001000111111010111111010110",
    308 => "11000011001000110101110110010100",
    309 => "00011111001001010011010011100000",
    310 => "00001101101011110101011001101100",
    311 => "01011001101001100011110000001010",
    312 => "10100001101110100010101101101000",
    313 => "00000101101100001000111110101010",
    314 => "11001110001100101011010110100100",
    315 => "10000111001101101001110101110110",
    316 => "10100111100101001110100110011010",
    317 => "00111100100100110101011110110100",
    318 => "10100001111000110100000011100110",
    319 => "01100000101010110110111011000010",
    320 => "00100110010110101101111100110010",
    321 => "00100100100010110010010111110000",
    322 => "10101111000000111001111001100010",
    323 => "10011011100100010100001110110110",
    324 => "00110100000101110010001001010100",
    325 => "10101110111001100000010101100000",
    326 => "11010000100000111000011011100010",
    327 => "01010111001001111011001001110010",
    328 => "00111011011101110011101101101110",
    329 => "00100000100011110110011001011010",
    330 => "01011111000010101000100111100100",
    331 => "11001100100001011111110111000110",
    332 => "00110011000001001010011101110110",
    333 => "00110111100010010010010000110110",
    334 => "01000101100001010001001010110010",
    335 => "11111011001101001111111111010010",
    336 => "11111101100111011100011101000110",
    337 => "11111000100110001101100100101100",
    338 => "11100000100101101101100111100000",
    339 => "10100001111011010010000001101110",
    340 => "11010010000100100101110110011000",
    341 => "01011001101001011011011110101110",
    342 => "11011100100010101011011111011010",
    343 => "10010111111110111100000001010110",
    344 => "10010000111101000100111110011110",
    345 => "10100100101111011100100100101110",
    346 => "01100011100000001011001001101100",
    347 => "11111001101011110000010011110110",
    348 => "11111101100001100011010101100110",
    349 => "01101110100000011001100101010110",
    350 => "11001100100101111000100101001010",
    351 => "10110010000001010000001101010110",
    352 => "10001100100110111011101111011010",
    353 => "11111010000010000011011000010010",
    354 => "01000001111101101111001011001010",
    355 => "10000101000100111101001101110010",
    356 => "01101111110111100100111010101010",
    357 => "10111001101011001101011111000110",
    358 => "10010010101111011110101111110000",
    359 => "01100111100010000101000101110010",
    360 => "00001101010001001110100011111110",
    361 => "00010110110001100011100100100110",
    362 => "00000000101011000011110100100010",
    363 => "00001010010100111110000001000110",
    364 => "11000100111011000100001010111100",
    365 => "01000100010100001111100111001000",
    366 => "01100101101000101011011111001110",
    367 => "01011110111010111111110010010100",
    368 => "00100100000100100101101110110000",
    369 => "01100010101001000101000011101000",
    370 => "01111000000001010001101101011000",
    371 => "01111101001000101110011100110000",
    372 => "11001001101000110111000100101010",
    373 => "00110111011011101101011010100010",
    374 => "00001011101001010001100100100100",
    375 => "00000011010000110110101110010100",
    376 => "00101110010110011001000001111100",
    377 => "00001100111000001001001100100010",
    378 => "10101101101111001101011101000000",
    379 => "00110000011100100011111111111010",
    380 => "00010011001001110010000010100000",
    381 => "00000111010100110011010000010100",
    382 => "01101110001100101101011110100000",
    383 => "01101110010000011001111111111000",
    384 => "11000010010010101111110100111110",
    385 => "11111011100000100011000010111110",
    386 => "00111011110110101101010001111100",
    387 => "00100101010010110100101111100100",
    388 => "00110010101000001111011000110110",
    389 => "11100101000110110001110101100000",
    390 => "01011010100000001000100001100110",
    391 => "10000101101000111110100001000000",
    392 => "01011111011001000111010110011010",
    393 => "00000001101011001111111000111010",
    394 => "10101001001111001011000111110000",
    395 => "10000111101011110111001110011010",
    396 => "10010000111001010100001011000000",
    397 => "10011010000010010011011011010010",
    398 => "10001011011011110000001010011100",
    399 => "01010011010000100001101000010110",
    400 => "10011001110000110011101100110000",
    401 => "00000010101000101000001011110010",
    402 => "10010111110100001111111001111000",
    403 => "00011111000001101001111101101110",
    404 => "01110110110000111110100000100000",
    405 => "11101000100010110111010011101000",
    406 => "11001110000111000001011001111100",
    407 => "10111011101100110000001001001110",
    408 => "10100100110000101010101101000010",
    409 => "11000000100001000001100100000000",
    410 => "11010101100001010011101001011110",
    411 => "00000001110011100101110100101110",
    412 => "01000001010001101101001011011100",
    413 => "11101000101011010101010100110100",
    414 => "01111011010011111001110010100000",
    415 => "01010110101101110101111001110000",
    416 => "01001110010001110100100110100100",
    417 => "11010111011001011010000010111010",
    418 => "10010001111000010010001101100010",
    419 => "11100110001110001101110101011110",
    420 => "00010111010101011000001110110010",
    421 => "11011101000100101110111100100000",
    422 => "11000000000111100011011100101100",
    423 => "10010110001000000000011011001100",
    424 => "01011001011011001000100010100000",
    425 => "00110110000111111000010010000110",
    426 => "00100010000001000101000100101000",
    427 => "00011000011101011011000001110100",
    428 => "01010111000000110010110011011110",
    429 => "10110011001000011110110011011000",
    430 => "11000000010000101011100000001010",
    431 => "01101010100101000001000000010100",
    432 => "01100110100000110110001100101110",
    433 => "01110111111001101110001001010110",
    434 => "00111011100010011001110010111000",
    435 => "10000100001001110110010001111100",
    436 => "10110000000101010101101000100110",
    437 => "00111011100001101101101001010000",
    438 => "11111101001100010100100101001010",
    439 => "01011000010010100101011001001100",
    440 => "10101011011101110010011100011100",
    441 => "00001000101001110100111011111110",
    442 => "01001001100101010011110000010110",
    443 => "00110011110101101001110000010000",
    444 => "00100101011010101010011101110010",
    445 => "11110110000010100100000011111110",
    446 => "11110100000100100011010110101000",
    447 => "11110111011111101011101110010100",
    448 => "00100101101100111011011000100110",
    449 => "11010110000011110110110110100100",
    450 => "11010000100111110100010100010000",
    451 => "00110111001111100111011010110000",
    452 => "00111110101000010110111000110100",
    453 => "01110100000110101101001000110010",
    454 => "11000111100100110001010001010100",
    455 => "00010101101001001000001101101110",
    456 => "11011110000011110001110100001010",
    457 => "01000011100100101000101110101100",
    458 => "01000010100110100110000001010100",
    459 => "11001011010110101001001110000000",
    460 => "11100001100101010110010010010100",
    461 => "11010000110111011010100000110000",
    462 => "00100101000111111010010101110010",
    463 => "10110011010110111111010100010000",
    464 => "00111010110010001111111001111010",
    465 => "00101111010000101111111010100110",
    466 => "01100110110010101011010000001000",
    467 => "00001111010101001110011111011100",
    468 => "01011100100001101100011110000110",
    469 => "01100100100010000100011000101110",
    470 => "11010011000100000100000010010000",
    471 => "00011010001101001100000001010110",
    472 => "10011011101010000101001011000100",
    473 => "11011011111011111100011000111100",
    474 => "11011000011010000001100111011000",
    475 => "01001001100001001100000001000110",
    476 => "01101011110010101110001111000000",
    477 => "00010010110001111101010010100110",
    478 => "11100101110011011110100010000000",
    479 => "01011111000001110011010110000100",
    480 => "11010010101101111010111111101110",
    481 => "10101111001101110010000000101010",
    482 => "11111000000010010110011010001010",
    483 => "01100010001010100000111100111000",
    484 => "01000101001011111100101000000110",
    485 => "01111011101101101000011100110100",
    486 => "11000100000011001100010010100110",
    487 => "11001100100011101010101000011010",
    488 => "01110111000000010010100011100110",
    489 => "11000001001010001001001001001010",
    490 => "01010010111010001000010100111010",
    491 => "10001100100001101001111111110100",
    492 => "10101000001001110100011000010010",
    493 => "01010010110100000111010101010110",
    494 => "01101000100111010100100100011010",
    495 => "00110001110001100101100111100010",
    496 => "01000011010000001101001001111000",
    497 => "11111000000110001001001010010000",
    498 => "00100010110001101001110010100100",
    499 => "10010011000000110000111000001100",
    500 => "10100100001000110101101000011000",
    501 => "00000011100000011000101010110010",
    502 => "00100111110110011110101111000100",
    503 => "01001011000101000110001010101010",
    504 => "11111011100111001100101101110010",
    505 => "11110001010011100010011101110000",
    506 => "10011010000101110110010011111000",
    507 => "10010000011010010111101111101100",
    508 => "10100000010000010000111001111000",
    509 => "11010011100000000101000011110110",
    510 => "00011000001100010000110010011100",
    511 => "11000111100000011001111111011000",
    512 => "11101001100000011010101010001100",
    513 => "10011010000000100101001000001100",
    514 => "10011101000010110110110110010010",
    515 => "11110111011111011101100011001000",
    516 => "00111110110010001111111001100110",
    517 => "00101100100011110001100010110000",
    518 => "11001110000100011101100000101100",
    519 => "10001000100111110111101110011000",
    520 => "00000111000100011001110000100110",
    521 => "10011011011001000011101000011010",
    522 => "11111011000000001001111011011110",
    523 => "11100110100110010100000010111110",
    524 => "00010010001001011111001101111110",
    525 => "00100111010010011001000110100010",
    526 => "01000010100000110011001100011110",
    527 => "10001001000100010100011110001010",
    528 => "10110001100001101110010010011000",
    529 => "00111011010101110101100100110010",
    530 => "01010011000110111011000100000100",
    531 => "00010010111000010010000101110110",
    532 => "00110000110110001001100000101100",
    533 => "01111011101110110101101111111000",
    534 => "00111010001100011011101110110000",
    535 => "01001011110000010010110001111000",
    536 => "10000001100011001100010111110100",
    537 => "01100101100110110110000111001010",
    538 => "00010110000110011011111111010110",
    539 => "00011010111000111000000010000010",
    540 => "10001001100000010001000001111010",
    541 => "01010101110101100000001000000000",
    542 => "00110100000111000001001000111100",
    543 => "11111011000010011001110110001110",
    544 => "10000101000101111111000101000010",
    545 => "00110111010010010100001111110100",
    546 => "01101100010011010110100100110010",
    547 => "11101101010011010100011110111110",
    548 => "00001100101111111011101110100010",
    549 => "10011111001110110111110000100010",
    550 => "01110000101000011000010000010010",
    551 => "00001011100000011010111100000010",
    552 => "11010101011000010000100100011100",
    553 => "01110001110100110010011101000110",
    554 => "01000000100000111111110010111110",
    555 => "10010110111111010110001011010110",
    556 => "11010010000100111011100101111000",
    557 => "10011001000010011100101111000010",
    558 => "11001110110110111100010000101110",
    559 => "11101111000001011111000010000110",
    560 => "11001101100100001101111010100100",
    561 => "00101111010110010010100100101110",
    562 => "11110011101000001100010100111100",
    563 => "01011010001100011001010010000010",
    564 => "10001000111101100100111000100010",
    565 => "11001010100101100101000100000000",
    566 => "11100111101010101110110100100000",
    567 => "11101110111110010001000000000000",
    568 => "11001010010001010001111011100010",
    569 => "00101011101100100000011110000100",
    570 => "11110000101000100011110111000110",
    571 => "11010111110111000110111000010100",
    572 => "10110010100110101011001100111010",
    573 => "11001100000110000000001011100100",
    574 => "10001000000100110101101110110000",
    575 => "11011000100110010101100011110010",
    576 => "01100100100011111110110111000010",
    577 => "10010010101010001010101110000100",
    578 => "10100111110010001110100110001100",
    579 => "11011011110001010010011000001000",
    580 => "11101001100100001110110101010010",
    581 => "00101101100001000001101000101110",
    582 => "00010001100001101100011010101010",
    583 => "11010111110100101001010101000110",
    584 => "10000011000011110101110010010010",
    585 => "00110110111010011101100001110010",
    586 => "10100011101101110101100111110110",
    587 => "10111010010010110010010010000110",
    588 => "11000001001110100100100110010010",
    589 => "00000100100111000100110100111000",
    590 => "00011110000011111111111000001010",
    591 => "10000001001001111111111001001010",
    592 => "10000111011001011001100111111110",
    593 => "11111001101110110111011001010000",
    594 => "00000110100011000101101001101000",
    595 => "01000101010111110111101100111100",
    596 => "11000110110010011011000110110000",
    597 => "01010011001011001111011101000100",
    598 => "10010111001110010011000001111000",
    599 => "00111011010010110101000011001000",
    600 => "01011101111011101010001001010100",
    601 => "11010011000111110010010110111000",
    602 => "01111000011000100000001010100010",
    603 => "00110000100111111100000001101110",
    604 => "00100011100011100101100110101010",
    605 => "01100010100110100011110001110010",
    606 => "01001111101101110110001011011010",
    607 => "10001010100111010011011111000010",
    608 => "01000011111111100111011000011110",
    609 => "11001011001101111101110110110000",
    610 => "00101110110001010101000001011010",
    611 => "11010011110000000001011111101110",
    612 => "01101010101000011011110110000110",
    613 => "00111111111101011011001110100110",
    614 => "11010101001010011011010100010100",
    615 => "10011111011000011110011111001100",
    616 => "01110000100110101011000100001100",
    617 => "00110111111100111100000001110100",
    618 => "10000011000111101111001101101000",
    619 => "10100101110001011100001000000110",
    620 => "00100001000001110011101010110000",
    621 => "11101011100000001111010001011010",
    622 => "01101111011000001111011001011010",
    623 => "01001011000011100011100101000010",
    624 => "11111101100111110100001010001110",
    625 => "00000001000000011010111100001100",
    626 => "00101010000100111111011101001110",
    627 => "00100101001011011111011111011000",
    628 => "10011001110010000100110110001010",
    629 => "01100011100011010001011000110000",
    630 => "10001010010100111011011000100100",
    631 => "10101110110111100000010000000010",
    632 => "01000000010010111010100100011110",
    633 => "00101110000001011110000011111010",
    634 => "01011011110110100101001010100010",
    635 => "01110001101010100000001000011100",
    636 => "11000010111010011111000001001100",
    637 => "11000000100100001000011100101010",
    638 => "10010111100011110011000101111100",
    639 => "00100111011010111001100110111110",
    640 => "11101101110001110111000101000110",
    641 => "11110000011011111001010000011100",
    642 => "01101001011000101001111111010000",
    643 => "11111011010010011100110110111100",
    644 => "01000110100011001111100100100010",
    645 => "10111111100011001011110100110010",
    646 => "10110110001001001110011011001100",
    647 => "00010110010001110100100101011000",
    648 => "10100011100100110111111000111010",
    649 => "01011111101111000001101011111010",
    650 => "10010110011111110111101111100100",
    651 => "01001001111100000010010100011100",
    652 => "00110101101010010111101000101000",
    653 => "01101010100000001001101010010110",
    654 => "11001011110100101000010110101000",
    655 => "01101000111100010111100111100000",
    656 => "11100110100001110010101110011100",
    657 => "01001111110011000000011111001100",
    658 => "01001011110000100110110100011000",
    659 => "11010110001100101101111001011100",
    660 => "00101101000111110101111011001110",
    661 => "11100110010111010001110010100100",
    662 => "00000111010100010111010000000100",
    663 => "01011101000000100001000101110100",
    664 => "01000100000111000010111001000000",
    665 => "10101101100010010010111000110000",
    666 => "10010001010101100001000100100000",
    667 => "10110111000100110101011100101100",
    668 => "10000101000100001010110011000100",
    669 => "10010111011111101100101100010100",
    670 => "10110110100011011100111010000000",
    671 => "10001101101011000110000010100110",
    672 => "01011100110101100111101101110100",
    673 => "01110000000101001001101001010010",
    674 => "00101011110010101010110100000000",
    675 => "00111110000110111101001000101010",
    676 => "01011111001101100101001000011000",
    677 => "10111111011110001111101101100110",
    678 => "00100100010011011111000101011100",
    679 => "00010100101000011001011100010100",
    680 => "11011100010000010010000110010010",
    681 => "11000110001010000000110101010000",
    682 => "00111100101110010010100011110010",
    683 => "10110111110100000111111110010100",
    684 => "00100010000000001011011100000110",
    685 => "00010101111000010000100111011000",
    686 => "01010010110001010100111110001010",
    687 => "01111000101010110110110100111100",
    688 => "00000100001110111110001100001010",
    689 => "01011011011111111010101111100000",
    690 => "10110010001110101101110010111000",
    691 => "10001100001010110011101101110000",
    692 => "01000001001100010010110100000000",
    693 => "01111011001101101100101111110100",
    694 => "11101011001010000111011010010110",
    695 => "01010001001000110000101011000010",
    696 => "01010101001100100110000110011110",
    697 => "00111000001110110101010100010100",
    698 => "00010111101111010000011100110100",
    699 => "11010111000000011111011010001000",
    700 => "11000010100011000001111111100100",
    701 => "10010101011000010001010110000000",
    702 => "00010011100100111111100010001100",
    703 => "01001000000111100111100101000100",
    704 => "11111010000010101001111011101000",
    705 => "01001011000101001111110111100010",
    706 => "01000000010010110000011111100110",
    707 => "11000001000000001001011000110110",
    708 => "00100110000100110110110001011110",
    709 => "01101010001101111010110110100110",
    710 => "01001111001110100000100111111110",
    711 => "01011011111010000111011000010110",
    712 => "11010101111100100001101111111010",
    713 => "00111001100111010010100101000110",
    714 => "10000111011100010000001010010000",
    715 => "10101010100100011110000110000100",
    716 => "00000000100101100000110110000000",
    717 => "11100010011111001001010011011000",
    718 => "01010001001010000001100101010000",
    719 => "00101111001001110111010110010000",
    720 => "11010001010011011000010001010000",
    721 => "01111010101000010101111000011110",
    722 => "01010100101011110101000100111010",
    723 => "00010110010100110010101001110110",
    724 => "01111011000000100000100111010000",
    725 => "10001111001100000011010101111100",
    726 => "10111111001000110001000000010110",
    727 => "01110001110111010111100101110110",
    728 => "10000010011110101000001111110010",
    729 => "10000101111101100110010010100110",
    730 => "00111111001110010000101001001100",
    731 => "11010111000000011011110010000110",
    732 => "11110011100101111101010101101000",
    733 => "01010111001001111100101100001110",
    734 => "11100111000111100111000110110100",
    735 => "10010011001000100010100111111110",
    736 => "10000011110001001011011101101100",
    737 => "01001101001110110010011010000100",
    738 => "01001100100100101110110001110110",
    739 => "01010110100000101011101000011010",
    740 => "11100111010101111100110111110100",
    741 => "10010100111100100111101011011000",
    742 => "11010100000000100100010010011010",
    743 => "00111110101110010000100011011010",
    744 => "10110101100000000011101001111000",
    745 => "01100011011011101111111000011110",
    746 => "01111000010100100111011010110110",
    747 => "10110111101011100011011001011010",
    748 => "01110110111110000100001110001010",
    749 => "00110011111001100101011111000000",
    750 => "00011000011100111110100001010100",
    751 => "10011001101010011011110001110110",
    752 => "11011000000010011111111100001000",
    753 => "11110111111001100001101111011010",
    754 => "01001101101011111100100110000000",
    755 => "01101111010000111010000111101110",
    756 => "00110111001011001100000001100000",
    757 => "11011110101101110000010010010010",
    758 => "10001110001000100111000000111110",
    759 => "11100100101100101000000010111010",
    760 => "11100101010101000111101100111000",
    761 => "10111011100000110001111111101000",
    762 => "10000101101001010011000101000010",
    763 => "01001100110000010110100111000110",
    764 => "00000101001101001010101010111100",
    765 => "01011101110100001000001101001110",
    766 => "01001010111000111000110110000100",
    767 => "10111101000011001101101001110110",
    768 => "11100001100111101100110101001000",
    769 => "11001010101000100100001111110110",
    770 => "00000110011111111100101100010000",
    771 => "01100111100101011001111111111110",
    772 => "01000001010011001011010011010010",
    773 => "11001100000001001010100001000110",
    774 => "01100111000001110100111001000000",
    775 => "10010110001101101111110111001010",
    776 => "11111100000010001111010000010010",
    777 => "00101101001010001010010010101000",
    778 => "11001000000100000110000010110000",
    779 => "10000001100000000000001011010100",
    780 => "01111101110010001000100110100110",
    781 => "11101110000110101000011101011000",
    782 => "01011010000000100110000010001110",
    783 => "01101110101110010100011011001100",
    784 => "01100011001101100101000011101010",
    785 => "11101110000110111011100000100010",
    786 => "01110110100010101011010011111000",
    787 => "00101010100001111001110111110000",
    788 => "00011111001011101100100101010000",
    789 => "10001010100001010010010010011100",
    790 => "00101010010110001011000110100000",
    791 => "01010101101100000010000011111110",
    792 => "01110101100110010000001111111010",
    793 => "10101011001011100011001010000100",
    794 => "10001110000111000111010001010000",
    795 => "10001111000101101101101011100010",
    796 => "01001001101010111010101111110100",
    797 => "00101010100100001101111110110100",
    798 => "00100111110011110001100011101010",
    799 => "11110101000010111011011010111100",
    800 => "11111010101000100110101100101110",
    801 => "11101110110011110100011110001100",
    802 => "10100110100100000100101111100100",
    803 => "00011110110001111100110000011010",
    804 => "10010111011100100101100000010010",
    805 => "11010100111110110101010000001000",
    806 => "01110010101010010010100111011010",
    807 => "01110011001011001101000111100010",
    808 => "00001011011000001111111111010100",
    809 => "01001101101100000100010000010010",
    810 => "11110100001110001111100000000100",
    811 => "10011000111011111110111110010010",
    812 => "11001001000011010111001001000100",
    813 => "01111001100100100111000001001000",
    814 => "01010100011111101010101111101010",
    815 => "10001010000001001110100011001000",
    816 => "01011101010010110110110111000010",
    817 => "01110111011101001110101111010100",
    818 => "10001010000010011001001000000100",
    819 => "10111000000101000000011011000000",
    820 => "01100010100011110001010000111000",
    821 => "00010001101100110110010000110000",
    822 => "11011010101100011101001011001000",
    823 => "11110110010001110010010111010110",
    824 => "01111011010101001101100011111100",
    825 => "00000010101111010110110011111100",
    826 => "10100100000001111010011100001110",
    827 => "10110000101011110001101010000010",
    828 => "11100010010011000110011111010010",
    829 => "11100001000100101101111001011010",
    830 => "00011100000011101111011011100110",
    831 => "10001001000010110011010001100110",
    832 => "01100111000010111101110100011010",
    833 => "10011001110100110110111011010110",
    834 => "10010101100111110010100100101100",
    835 => "01001000101001000011001101110110",
    836 => "01010100110001001000100101001100",
    837 => "10101111100000111011001010101100",
    838 => "10001100101000100110110011101010",
    839 => "00010010010000010001010011100000",
    840 => "00011101100100111011000100100100",
    841 => "10101110001111100011001010100100",
    842 => "00100110100001100000011001111000",
    843 => "11111011101101100010010001101110",
    844 => "01001010100010011110111000110100",
    845 => "01110101110000011001100100111010",
    846 => "10010100010011011001010110100000",
    847 => "11010111001000100001100101101000",
    848 => "11010001000010101101011000011000",
    849 => "01010000011000001111100011101110",
    850 => "01110000100011110000001011010000",
    851 => "00010001001011000001000001101100",
    852 => "00111111100101101111100011011100",
    853 => "10010011100110000101001000001000",
    854 => "11101110101000100011010010110100",
    855 => "01011110110101010111001100011000",
    856 => "11011111010100011110100011011110",
    857 => "11011101101010011110001001011110",
    858 => "00100000110111111101011000011100",
    859 => "10010000100011111001100000011000",
    860 => "11110100011001101110111010010010",
    861 => "01000010000101110000111010000110",
    862 => "11100110010010111000011110000100",
    863 => "10100000100110000101001010001100",
    864 => "00001101011100001001010111001010",
    865 => "10100001001001001011101101111100",
    866 => "10001101001010001110101010010000",
    867 => "01000110100000110111111111011110",
    868 => "01110110001011011011101111111100",
    869 => "10011100001011001001111101001010",
    870 => "00000011000111001010110001001110",
    871 => "11110100001110111100011001100010",
    872 => "00001011010100001000011010000100",
    873 => "01101011100000010001010101110100",
    874 => "00101110100011111001101101011000",
    875 => "10011010101110101011011101111010",
    876 => "10000101100010001101000010110100",
    877 => "00101110110011011010000000111000",
    878 => "11111001001111110001001011101100",
    879 => "00100110010100000000010101101100",
    880 => "11000011100100101100010111110100",
    881 => "00000111110010110111111011011000",
    882 => "11111101000011000010011111111100",
    883 => "00100000101011100000100101101110",
    884 => "00101011100010111011100001011110",
    885 => "11011011001111010110000001101010",
    886 => "10111011000111000111001100000010",
    887 => "10010100010000011111100110011010",
    888 => "00100100101000010111100110111000",
    889 => "01110101110011110011101011101100",
    890 => "11111001010010110100110011001110",
    891 => "01110000100110010001011110110000",
    892 => "11110011011011110111011010110000",
    893 => "01111010101100110000101011101110",
    894 => "01110011101101001100111100111000",
    895 => "01100100011011000001010001100110",
    896 => "00010010001100101000110110101000",
    897 => "01001101000010000100010001110100",
    898 => "01010111110100110110011011110000",
    899 => "11110011000010011011101111011100",
    900 => "00101010010110010111101110111100",
    901 => "00000101110010000101001111111000",
    902 => "11110111101111000110000101100010",
    903 => "01000001100011100011110001101010",
    904 => "10000000110011111110100010011100",
    905 => "10000001010101010011010110100000",
    906 => "11001000000011011000010101101110",
    907 => "10100101100000000101011001111110",
    908 => "01011111000001111101000101100100",
    909 => "11011000010110010110000011001100",
    910 => "11100001101000000010010010000000",
    911 => "11010001100000011010010110000010",
    912 => "10100001010110100100000000010000",
    913 => "00101010000001000010100101110100",
    914 => "00011010001000111010101011000000",
    915 => "00101111100000111000000101001000",
    916 => "01001110010001100101100110101000",
    917 => "10000110010011101100010000101010",
    918 => "01100010111010110101000111000010",
    919 => "10110110110011011100111000110010",
    920 => "10001011100001100100001010110010",
    921 => "01100001000011010111010100110100",
    922 => "00101101010000100100111101111100",
    923 => "00010010001000001010001111000000",
    924 => "10101001110100000100101110100100",
    925 => "01100010001010100101000011111000",
    926 => "00101010011101111011110011010000",
    927 => "10000010100010011010001111110100",
    928 => "01010101010000000101100000110010",
    929 => "11001000001000001111101101000000",
    930 => "01001100101000001011111000000010",
    931 => "00110111000111000111001000011100",
    932 => "10110000000100010101001111011000",
    933 => "01100100001001110000001000100010",
    934 => "00001000100001011101110011110110",
    935 => "11111001110110110001000000001110",
    936 => "01010110010100011001101100001100",
    937 => "01101010101001101100110000001100",
    938 => "01100100100011111001100000011000",
    939 => "10010011000100110000011011110010",
    940 => "01101010100001101100000110010000",
    941 => "10011101000010110010110010000110",
    942 => "00101100000101001010101100111100",
    943 => "01100011111000001010111000011110",
    944 => "01001111001010110001011101001100",
    945 => "11110100000000110110101011100100",
    946 => "10100110110010100001111001100100",
    947 => "10111010000000011100111010111100",
    948 => "01101011101011110111110010000000",
    949 => "01101101000010000101100100110110",
    950 => "00111100010001111011100110111110",
    951 => "10001011010101110001000000111000",
    952 => "11000100111110011110000011011000",
    953 => "10011001011101011011001101000010",
    954 => "11110110000010100001110010001110",
    955 => "00111011000011001011101000001110",
    956 => "00100100111110010010111011110000",
    957 => "11111000100101111100110111100010",
    958 => "01111010101111001000011011100000",
    959 => "01010101100011100000110010000000",
    960 => "00001011101001001001010111100010",
    961 => "11101001000000111100000000010110",
    962 => "01110111101111111101010000000010",
    963 => "00001100100010100101111001110010",
    964 => "11000100001101000100000010110110",
    965 => "01011010110110111101010001111100",
    966 => "01100011100100000101001000100110",
    967 => "10010110010101000110111011001110",
    968 => "11011111011011010000011111010100",
    969 => "11010101000111110111000001111100",
    970 => "01011111011110001000010011101000",
    971 => "10111001000101111100000111010110",
    972 => "01101011011011000101000000111000",
    973 => "11011000100011011011000010011110",
    974 => "00010001010101010111111111000010",
    975 => "00110011010001011010000000001110",
    976 => "01111010101111000101101001111110",
    977 => "11010010101000100110001010100110",
    978 => "01000010010111011110011010000000",
    979 => "11011001001011000010100001110100",
    980 => "01011011110111011100011111110110",
    981 => "00001010010010001010010100010110",
    982 => "10011101011111100101110110001110",
    983 => "01101011000101000100100000101010",
    984 => "11010011100101000010011001011110",
    985 => "01010101011110101111011101000010",
    986 => "11010011100100011011011110111000",
    987 => "10111010100011010000000100111110",
    988 => "11000011011011001111101101000000",
    989 => "00101000010001111100101010110000",
    990 => "11000100010011111110101010111010",
    991 => "01110100111101111010000010000010",
    992 => "01111011000011010000100010101110",
    993 => "00110100110001110101110100110110",
    994 => "10101001111101101110000111000010",
    995 => "11000111001001011111000001011010",
    996 => "11000101001100111111001010111000",
    997 => "11001000011001001011010010101110",
    998 => "11110101010001001111101111110100",
    999 => "11100010101010001110101101101110");


  component finv is
    port (A : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          Q : out std_logic_vector (31 downto 0));
  end component finv;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (3 downto 0) of std_logic_vector (31 downto 0);
  signal cc : std_logic_vector (31 downto 0) := (others => '0');  
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0'); 
  signal Q_buff : std_logic_vector (7 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
  signal i_isRunning : std_logic := 'U';
  signal i_result : std_logic := '1';
begin  -- architecture finv_tb

  i_finv : finv port map (s_a,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk,Q_buff) is
    variable ss : character;
    variable count : integer := 1;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      s_a <= a_lut (addr);
      cc <= ans_lut (addr);
      ccc <= cc ;

      if i_isRunning = '1' then  -- rising clock edge
        if ccc = c and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 1 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;

  end process ram_loop;

end architecture;
