library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity floor_tb is  
  port (
    clk : in std_logic;
    Q : out std_logic_vector (7 downto 0));
end entity floor_tb;

architecture testbench of floor_tb is

  type lut is array ( 0 to 999) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "11111011101111011110001101010010",
    1 => "01110111111011111000000000001111",
    2 => "01111011110111100101111001000011",
    3 => "11011101100111011001011110100100",
    4 => "11111101001101111110101111101000",
    5 => "01111111011101101101100000001101",
    6 => "10111111111011111001010111100010",
    7 => "01101111011110101010111110111111",
    8 => "01011110110101100101110010001011",
    9 => "11011010011111101011100010010100",
    10 => "11010011011111101111010011111111",
    11 => "11110111010111001100010101001010",
    12 => "10110110111111010110111010101110",
    13 => "11111100111110111000001001110001",
    14 => "11011110101110111001101011101111",
    15 => "01111111010111011111101001001011",
    16 => "01111011010111111001100111100110",
    17 => "11111011101010101111000100101100",
    18 => "10111011111100101011001100101001",
    19 => "10101010110001011000010011100101",
    20 => "10110111011011100011011001101111",
    21 => "11011110111110110111110100011111",
    22 => "11111011111011110010010101101000",
    23 => "11101110111100101111100011010110",
    24 => "01101111110101011101000000010110",
    25 => "01110110111110111010000100100011",
    26 => "01111111000111110010001111111111",
    27 => "01111110111111111111000100110001",
    28 => "11101111011111111011101001010100",
    29 => "10111111110110101001100010100110",
    30 => "01010011111101010011010001010000",
    31 => "10111101011101111110101011100001",
    32 => "11110000111110001111110010110101",
    33 => "01110111101011001101001111111101",
    34 => "01010001010111111000010110101111",
    35 => "10101111111111111100011000011110",
    36 => "11111011100111101000011011010000",
    37 => "01110110111111101101011000111000",
    38 => "01101011001011111010010011011010",
    39 => "10010111111010111011001101101110",
    40 => "01101101110011100010100101110101",
    41 => "11011010000111110010000100100010",
    42 => "11100100111001000001100101000010",
    43 => "01011101111101110000110111101010",
    44 => "11111010111110111111100001011001",
    45 => "11111101011111100000011011001001",
    46 => "11111010111111111101100100110100",
    47 => "11111111010101010010101111100011",
    48 => "11110011111101011110100001011000",
    49 => "10110010100100010011001001011010",
    50 => "01011011101111111011110011100110",
    51 => "01101111111010110010011101101100",
    52 => "11011011110110110010010010101111",
    53 => "01001110111101001111011111001011",
    54 => "01101001111100110001000000111111",
    55 => "10111101111111111010111101110011",
    56 => "10110110011111110001011011110101",
    57 => "11110111101110111010101010111001",
    58 => "11111110111011001001000100000010",
    59 => "11111110111001110100111100001100",
    60 => "10011111000111110110111110011010",
    61 => "10100101111111101010000111111000",
    62 => "01011111111111110100101100100110",
    63 => "01111010100100111011101101111001",
    64 => "11111000011111111100000010011110",
    65 => "10111011111011110100110101101101",
    66 => "10111111100011110010111001001100",
    67 => "10111111111010011111011111101011",
    68 => "11100111110111100101110010110101",
    69 => "01110011111010100100010001010011",
    70 => "11111110111111000110001111010011",
    71 => "10110110110111111100000111111000",
    72 => "11110011011101011010101110000010",
    73 => "11011100111111100001111001001011",
    74 => "01111001011100011011110100010001",
    75 => "01111101101111101110101100011010",
    76 => "10111011111110111101110000000011",
    77 => "01111111011101010101100010110011",
    78 => "10110111111111110110010000100010",
    79 => "01110111111111011011111101111100",
    80 => "10110111111001111100010110001011",
    81 => "01110010110001001100010000100010",
    82 => "01011011011101010101111011000101",
    83 => "10111101111111111001010111101010",
    84 => "11111011111111111111011110000001",
    85 => "11111011111110011010101011111011",
    86 => "01011110011111101010110010011100",
    87 => "10111111110111110011110010101110",
    88 => "01111010111110110111000110011010",
    89 => "00111111111010110010001100011011",
    90 => "11100110111111101010011100110110",
    91 => "01011111100101011100100111011111",
    92 => "11101101010110111000011011101000",
    93 => "01101100011111110101001110001011",
    94 => "10111111101101110110111010110011",
    95 => "01011111101010110101101111100110",
    96 => "01000110111111011111111001011010",
    97 => "11111110111101111101000100011100",
    98 => "01001111110010110101110101011111",
    99 => "11111110111111110100000111010110",
    100 => "10101100111110110111001100100111",
    101 => "10011111011110111010010011000100",
    102 => "01101111101111010100101100101000",
    103 => "10111110111100110010000011010110",
    104 => "01111011100110100111100000100000",
    105 => "11100111110111001011011001100000",
    106 => "11010110111010110000000100011111",
    107 => "01111101001001011110101101110001",
    108 => "11111101111011101110111000100101",
    109 => "10111111010110110110001111100111",
    110 => "11010111010111101001010011000010",
    111 => "11110110100111001100110100001011",
    112 => "01110111111011111001000001000000",
    113 => "11011111111111100011101110001010",
    114 => "11101110111100110110001011111110",
    115 => "01110010110111110011001011000001",
    116 => "11110111101111111101101111001000",
    117 => "11101100111011000000001100110011",
    118 => "01111110101000110100101010000101",
    119 => "01101111101111110101001010000101",
    120 => "01000110101110101010100010101010",
    121 => "01011111100101010011011101100101",
    122 => "11111100101101111111111111101011",
    123 => "11011100111111101100110111010111",
    124 => "01111110101110011010001011000000",
    125 => "11011110110010100000001011000110",
    126 => "01101101111001111110101111111110",
    127 => "01011110101111111000110011111011",
    128 => "01111011110000111001011001011110",
    129 => "01011110111111001111011001000101",
    130 => "11111011011110011000111110110011",
    131 => "10110011111001110111010011001100",
    132 => "11010110111101111101000101011001",
    133 => "01101011111111101101110110001010",
    134 => "11001111101101100010010010001100",
    135 => "01111011111110010110010010001000",
    136 => "01111101011111111001001011000101",
    137 => "01100111111111110010100000011001",
    138 => "11111011111110110011000101101010",
    139 => "10101111101101111010100100100011",
    140 => "10111111101111011001111011100010",
    141 => "01101110101101111000111011000111",
    142 => "11111110011010111011100100110000",
    143 => "01101101111111101000001111101100",
    144 => "01010101111011010110100000001110",
    145 => "01010101111111110000010011110000",
    146 => "11101101100011110100001000100000",
    147 => "00111111110010111010011110111010",
    148 => "01000101101111110010100010010111",
    149 => "11110110100010100101011110100001",
    150 => "01011001111011111011000111000010",
    151 => "10101001001001011101011011101111",
    152 => "01111110111111111001100011101111",
    153 => "11011111110111111111111001001010",
    154 => "01110111111111111000010010010110",
    155 => "01110001111111111100011101011011",
    156 => "01011100110111010101010100011011",
    157 => "11010111011111111010111011110101",
    158 => "01111111001101111111101001010000",
    159 => "01111011101100010000101011000101",
    160 => "11111011111111111110110000001001",
    161 => "11101111110101011111010000101101",
    162 => "01101111001011110000011010101011",
    163 => "11111011011111011110001001011000",
    164 => "10111101011111111011000001110110",
    165 => "11101110111001010111110011100010",
    166 => "01001011111111010101101000101101",
    167 => "01100011111010110010011000101111",
    168 => "01111001101100110001001010000101",
    169 => "01011111010010100110111011110101",
    170 => "01011010111111111101101101010011",
    171 => "01101111110111111100111111001001",
    172 => "11010111111101110110111110100000",
    173 => "01110110010110110101101101011100",
    174 => "10011011001110010010111010111000",
    175 => "01010110111101110100010100100110",
    176 => "01111011111111110000111001100110",
    177 => "01101010101111111010010001011101",
    178 => "11101011101111010100110101010111",
    179 => "10011111011110111000101000011100",
    180 => "11111011111111110100010111010111",
    181 => "01111110010111011010000000000011",
    182 => "01111101111001010111010110100111",
    183 => "01001101011110110110100111110111",
    184 => "11011111100111111010101111101100",
    185 => "01110111101011110100111111100010",
    186 => "01111110100111110100010011111101",
    187 => "11101110011111111100010010100100",
    188 => "10010011111101111101000010110010",
    189 => "11111111001110010111111110111111",
    190 => "01111110110110010100011110101011",
    191 => "11010001110110101110111010101010",
    192 => "01111111010011111100101000110111",
    193 => "01101011111010111000110011011110",
    194 => "11110110111111100110011110101110",
    195 => "01110011100110110100011111110111",
    196 => "01111111010111101011111010010110",
    197 => "01111111011110010001101011100011",
    198 => "01001011101011101000110100010011",
    199 => "11101111100011001000110111100000",
    200 => "01111100100011101110100110001011",
    201 => "10111111101101100101011001010000",
    202 => "10011111111011010100101111010000",
    203 => "10110111011111110100000001110000",
    204 => "10011011111001111000000110101010",
    205 => "01001011010000011100011100011010",
    206 => "11101001111111111101100111000101",
    207 => "11111011110011110100000111011110",
    208 => "01101011111001111010100000111110",
    209 => "11010101011011100011100110010001",
    210 => "01111011110011010100001000100000",
    211 => "01101011111010111111101011110110",
    212 => "01010111111111111010000000001110",
    213 => "01010001011110111110000101000010",
    214 => "11011111111101101001111110010011",
    215 => "01110111111000000110000101111110",
    216 => "11110010101101110001101000110101",
    217 => "01111101010110111001000001010000",
    218 => "11110101100101101000011111110101",
    219 => "01011101111110011011110111111100",
    220 => "11100111101011110010101111001000",
    221 => "01111101101010101000100000111111",
    222 => "11111010000111100011001001000110",
    223 => "11110001111110100000111111110001",
    224 => "10101111101001001011011110101101",
    225 => "01111101111111111001000010111110",
    226 => "11101110110111111101000011000010",
    227 => "01110111010110010110000100000011",
    228 => "01111011111111100001101000111010",
    229 => "10101011100110101110001001110111",
    230 => "01111110011110101101011101001100",
    231 => "01011111011010111110001100011000",
    232 => "10100101011101100011010000001110",
    233 => "01111000110111100111110011011010",
    234 => "10111111111110001010000100110001",
    235 => "11001111111111101010011100001000",
    236 => "01101111011010111001111100100101",
    237 => "11111011111110111101101000000100",
    238 => "11111011111111100010100101010110",
    239 => "11110001110100111001001010110110",
    240 => "01101111111101111001100101111010",
    241 => "01101111001111110000100111001110",
    242 => "01101011111111010000110000001110",
    243 => "01111110111100111110011000001001",
    244 => "11111101010101011101000011010010",
    245 => "10111011111010101110110101101101",
    246 => "01111011111111110001110010010110",
    247 => "11011111011101110101010011111110",
    248 => "11111110011110011001000110001011",
    249 => "11111110111011101100001100101010",
    250 => "11111111001011110110011111011100",
    251 => "10010011111101101100011111111010",
    252 => "01011010111111001000011100100100",
    253 => "01110111101111110111001000110101",
    254 => "01111100101011110111111000100100",
    255 => "10001010101110101000101011011011",
    256 => "11011101111111111011000001111010",
    257 => "11101101010111001010011001001011",
    258 => "10010011111110111000101000110011",
    259 => "11101111110011010011010100110110",
    260 => "10101111101101011011010100110100",
    261 => "01111110111100010100000000111010",
    262 => "11010111111001011000000001100101",
    263 => "01000111110111110111111101010100",
    264 => "11110111001111111000111000110010",
    265 => "01010111011011111110000010111101",
    266 => "01110111111111110111100001100010",
    267 => "11101110100111111011000011011100",
    268 => "01111111001101011000100010000001",
    269 => "01110011110111110110011010011010",
    270 => "01111101111111101011100100110011",
    271 => "01111101101011110011101010110100",
    272 => "11111001001001110001101001001011",
    273 => "11111101111111101110101011111010",
    274 => "01111101111111010100101101001000",
    275 => "10101111110001111010101001100110",
    276 => "11110101110110010010001100100110",
    277 => "01111111001101111101011100110001",
    278 => "11111100111111111011011011111001",
    279 => "11111101110011111110011101100011",
    280 => "11101101111101110101001011010111",
    281 => "10111101100010111110111000110010",
    282 => "01011010111111100000101001000100",
    283 => "11110101001111110110111010001011",
    284 => "11111111011011111010110011111100",
    285 => "11111000011011100001010101110000",
    286 => "10111111111101100000110100110010",
    287 => "11110111111111111110101010100001",
    288 => "01111110111111110110110111100001",
    289 => "01000111110111110101100001000110",
    290 => "01011111111011011010100000010010",
    291 => "11011110111100000001100000101110",
    292 => "11111111011111010110111110010101",
    293 => "01011101111001111010000000100111",
    294 => "10111111111011110111111011101001",
    295 => "11101101111111010110011001000101",
    296 => "11011101111010110000101110000110",
    297 => "11101111011111010111010011110001",
    298 => "01011111100111100101101111001010",
    299 => "11011011111111110011011000111011",
    300 => "10111111110101111011100010001101",
    301 => "01111110110111110000111010111110",
    302 => "10110111111001101110111001001101",
    303 => "01101110111110111011111110101011",
    304 => "01011110101110110111001000110100",
    305 => "11101101111110110000011000001100",
    306 => "11100110011111000100111110001111",
    307 => "11111110111111010011111110010001",
    308 => "10111111111111100101000010100000",
    309 => "11111000111010111011101111101101",
    310 => "11010101100111111010010101100110",
    311 => "11111110110110110101001111101100",
    312 => "10101010111011110111100111101001",
    313 => "10111110110111010001100010101001",
    314 => "01110110111101101001001100010101",
    315 => "01111011111100010100001000101001",
    316 => "10110100110111110000110101110010",
    317 => "11010111101110011011100110110010",
    318 => "11111010111110110111101110001110",
    319 => "11110100010011110001011110001110",
    320 => "10110010001111111111100101000110",
    321 => "01011101111111101011101001011010",
    322 => "11111110100101110110011010111001",
    323 => "11111001111011110111011101000110",
    324 => "10111001111111111111011011111001",
    325 => "01110100111110110100110010010000",
    326 => "11111001101111101111111000000101",
    327 => "11011101101011111101100110101100",
    328 => "01110111011111101101101111101111",
    329 => "11110111100011000101011111101000",
    330 => "01101111011111101000100111100001",
    331 => "11010111011101110111011010010000",
    332 => "10110111101101110110010100101110",
    333 => "11011011111101110001001010010001",
    334 => "11001101110111001001011110110111",
    335 => "11101110101111101100010110110110",
    336 => "11111111000101111001001100011100",
    337 => "11111111011001110000111111001001",
    338 => "11001111101101110111110010100010",
    339 => "01101111111111110010111100011110",
    340 => "10111111101011101010001000101110",
    341 => "11111011110111111111000011111000",
    342 => "11001111111110101101011010011000",
    343 => "01111011110011101100110111010100",
    344 => "11110011011011110110100100000110",
    345 => "11111101111111000110101000111101",
    346 => "10111101110001111000111101101101",
    347 => "01110010111011111101111110101011",
    348 => "11111111011111100101111010011001",
    349 => "01001011111110111111110101000011",
    350 => "11011001001110111010001001010110",
    351 => "10011111111101111010001011000011",
    352 => "11111011111001110000101011001011",
    353 => "11111101111110011111010000010110",
    354 => "11111101100011100111011110001111",
    355 => "01001110101111010100000010111101",
    356 => "01001111111001111000100111101110",
    357 => "10111101100111001110111011110111",
    358 => "01111111001101010001000000100011",
    359 => "11011111110111000101111100000001",
    360 => "01111110111011110000011010111001",
    361 => "01100101111110111100001000011010",
    362 => "11011111101111110010111000100000",
    363 => "01111111011011110111100011110101",
    364 => "01011111011010111101100111011011",
    365 => "01111100101111110000001101110111",
    366 => "11010111111111110100111010000000",
    367 => "11101111011110001011101100111011",
    368 => "01110011000101010001010000111000",
    369 => "11111110011101100000101010001010",
    370 => "11111011110100110011000001111011",
    371 => "11011110111001000101001010110110",
    372 => "10100010110011011100110101110000",
    373 => "01001011111111010010011011110100",
    374 => "01101011011110110101001100000011",
    375 => "11111110111101011000100001101100",
    376 => "11111110111111110011100010101101",
    377 => "11110011111011111000101000111011",
    378 => "01101100111111001001110011111101",
    379 => "10110001101111011110111111100010",
    380 => "11111111011011010010011000000101",
    381 => "01011110100010000100111101011011",
    382 => "01100111111111001001011100011110",
    383 => "01110111111011010000110111100010",
    384 => "11011011011100111010000000010011",
    385 => "01011110111101100001100110010101",
    386 => "01011011110011111101011011100011",
    387 => "01100000111110101101111000100100",
    388 => "01101100111111111011011010101110",
    389 => "01111011111011110101010011011001",
    390 => "01001111101111110110110101001111",
    391 => "10111111111101000000010011100000",
    392 => "01011100111110110011111100101000",
    393 => "11101010111100101101001101011010",
    394 => "11110011011111110111100110111010",
    395 => "01011011111011011111100000111111",
    396 => "01010011110111101011110010001111",
    397 => "10110011011110110111100010100011",
    398 => "10111110111011111001000101001001",
    399 => "11111011110111011111100011000001",
    400 => "11110110111101111001010001110000",
    401 => "01001111001111110001101001111101",
    402 => "01101111110111100011111101000101",
    403 => "11101100110111011001111011001001",
    404 => "10110111111110011011010000010010",
    405 => "11110011011110100011111111101001",
    406 => "11001011101111110010011001010000",
    407 => "10100010101110101010101010110000",
    408 => "10110010111111111010110001111011",
    409 => "01111011100011111011100111010111",
    410 => "01111011011110111011010011000011",
    411 => "01111010011111111111110001111100",
    412 => "11001111111001110100000110101100",
    413 => "01011011001111110100011101010010",
    414 => "01110001111111110001000101010011",
    415 => "01111011100111011010011001011101",
    416 => "01100111101111101101000100100110",
    417 => "10100101011111111111110100101110",
    418 => "00111111111101111110100011010000",
    419 => "11111000111111110111100001110010",
    420 => "10011110110101110110011011010101",
    421 => "01010011100101111010101111110100",
    422 => "01111001111111110011111011001100",
    423 => "11111110111101111011010001110101",
    424 => "01111011111111111100000101111010",
    425 => "11111101111101100010101100011110",
    426 => "01111101110010100111101101010111",
    427 => "01001010001001110100101110111100",
    428 => "11010011110111111010011100111000",
    429 => "10111100101011111001110101100100",
    430 => "01111011110110011111010011011110",
    431 => "11010111101001110000100100100100",
    432 => "01111011111111110100101100111100",
    433 => "11010011111011110100001101101010",
    434 => "11111011001111110101001001101100",
    435 => "10110011001111001011101111000101",
    436 => "01111000001111110101011011010000",
    437 => "01011111011111101001100111100000",
    438 => "11111100111111101101100101110100",
    439 => "01111100110010111101011001000000",
    440 => "11111101011000111001011011110001",
    441 => "01111101111111111011010100001100",
    442 => "11101001111110111001000110001100",
    443 => "10011011101101110111100000010110",
    444 => "01100111111111110110111111101111",
    445 => "10111111101010111010000100000011",
    446 => "11111100011111010111001010110101",
    447 => "11110111111010110111111011011010",
    448 => "11100001011110111000111010101101",
    449 => "01001010011100111100001110000010",
    450 => "11011111101000110011001010011100",
    451 => "01111101111111011011010000110011",
    452 => "01111111010011011000100111010000",
    453 => "11111101101111110001100001101101",
    454 => "10111111111100010010110101000110",
    455 => "01101011110111110001010100001111",
    456 => "11010111110101110111011011111101",
    457 => "01110111110011011011001111111101",
    458 => "10011101011101111100010111001100",
    459 => "10111110101110110111111001101001",
    460 => "10101111010010111010100010010001",
    461 => "10011101111001000010111010010111",
    462 => "11110010110111101000100100101000",
    463 => "01110110111110110001001001111100",
    464 => "11101101111001101110010001011010",
    465 => "10000111001111101101110001010101",
    466 => "01010101011101111111010101100110",
    467 => "01011110011111011010111011000011",
    468 => "01101101111010010110101000010001",
    469 => "01110110000110110101011101101011",
    470 => "10111000111110011110101101101011",
    471 => "11011111111111111100101111110001",
    472 => "11111110101111010100101000111100",
    473 => "11110011011011000010100010111100",
    474 => "00111111111110011101110101010011",
    475 => "11111111011111111110011001011101",
    476 => "11110011100111110110011000100010",
    477 => "01111010111111010010100011000001",
    478 => "10111111111111111100110010110100",
    479 => "01111111011111110100011010001001",
    480 => "10111011101111101011010010010010",
    481 => "01010110100111111010000100111000",
    482 => "11111001101110110101110110011101",
    483 => "11110011101111011010110010100110",
    484 => "10011000110100110001010111011011",
    485 => "11100111110011010010000100100101",
    486 => "01101011011111110010110000001101",
    487 => "01010100110011111101110001010110",
    488 => "10111111111111110011111011000110",
    489 => "01110101001100111001000000000011",
    490 => "11111111011111011010011000010000",
    491 => "11101110111111110001100000110111",
    492 => "11101110111111100100000010100010",
    493 => "01001101111111111101001111101000",
    494 => "01011011111110110111011100001011",
    495 => "01111011101111111000100011001110",
    496 => "01111111001011111100101100001011",
    497 => "11111011111111101100011011110011",
    498 => "11111011100000110001101001010010",
    499 => "11110110111110100011010101011100",
    500 => "01111110011001110100011111001011",
    501 => "11110111110111111011000001010001",
    502 => "01110111011111101001100101000101",
    503 => "10110101011111011100110111110011",
    504 => "11111101110111110111111001101010",
    505 => "11110111111111010001101111101100",
    506 => "11111110101110110010000100010011",
    507 => "10111011010011111100111011000000",
    508 => "11110111011011110000011101000000",
    509 => "10111110011111111101001000110000",
    510 => "10111111101001100010100111101110",
    511 => "01001101010000010111101000010000",
    512 => "11101111111111001000110000100101",
    513 => "11011111111100000011101011101000",
    514 => "11101111011111100010001110001110",
    515 => "01111101111110010100000110011100",
    516 => "01110111111111110110111001001111",
    517 => "11101100111111111000100001000111",
    518 => "10111111111101110101111111101011",
    519 => "01111011011111111110001000101111",
    520 => "01001011110010110100100011101101",
    521 => "01111011110010010000100100010110",
    522 => "10010111011111010001000111100101",
    523 => "11011110100111110111011101000101",
    524 => "10110110011011100011001011100001",
    525 => "01011111011011110111000111111010",
    526 => "11011111011111110001001101000010",
    527 => "10110011101101111001011101101010",
    528 => "00111111101100110100010111010011",
    529 => "11101111111111110110111001001100",
    530 => "01011000011111111100001111100100",
    531 => "01101011011001110101001110111110",
    532 => "11111011111011110010010001111110",
    533 => "11011111111111110111001100010000",
    534 => "11010111110111110101000101110000",
    535 => "10010100111100100010001100000000",
    536 => "10010111111111111000101000001101",
    537 => "01111111011101111101101011000001",
    538 => "11101110111001001011001010110011",
    539 => "01101011100111010000011001111001",
    540 => "01001100110011010110111110010110",
    541 => "11011111111101110110100111001110",
    542 => "11010110000110110011101010000011",
    543 => "01111111001110110111011010000110",
    544 => "11111111011111111000110010010110",
    545 => "11101101111111110000100100010111",
    546 => "01011010111011110111010001110001",
    547 => "10110111111110011100010100001110",
    548 => "10111001111110110010110001101100",
    549 => "01111111000010111010011110011111",
    550 => "01111111011101110010100100111101",
    551 => "11011011101011001100100101010110",
    552 => "11111011111010011111010100010111",
    553 => "00111111111011111010010110010000",
    554 => "11110110110110010111100001000100",
    555 => "11011111011111110001000101110101",
    556 => "11011101111111111101010000001001",
    557 => "11011111100111111101101111100011",
    558 => "10111111111111110001110101011000",
    559 => "01011001110101101110100000110011",
    560 => "01011111110011110111010001010111",
    561 => "00111111111101100010100011100100",
    562 => "01010011011111101101101111001101",
    563 => "11100101011000110011001100101011",
    564 => "01101110111011111110010100101110",
    565 => "01110111101001110100101110110111",
    566 => "11111101111011111010000100101110",
    567 => "11111011111100100110010001001110",
    568 => "11111110110110110001001101000001",
    569 => "01101111101111111110001001001011",
    570 => "10110110011111100101110111101110",
    571 => "01111011111100011010101010011101",
    572 => "01111000111111010001000110111010",
    573 => "00111111110111111001011001100010",
    574 => "01110111001111111000010011011100",
    575 => "10111101001001111000110011000000",
    576 => "10111101111010011001111011111100",
    577 => "10011111110001111101111111011110",
    578 => "01111101111011010101010101000000",
    579 => "10111111101011110111011110011110",
    580 => "01111111001011011100011111010011",
    581 => "11011001100011011101010000100110",
    582 => "01111110111110011101010100010001",
    583 => "01111001111111010001010000101100",
    584 => "10101010111011001101110010111000",
    585 => "11110101110010110001000111110101",
    586 => "11111011001111110001001011011011",
    587 => "01101011101111110110101111100001",
    588 => "10111101111110110000111000101001",
    589 => "11101111010011110110110000010001",
    590 => "11000101110111100010111100000010",
    591 => "01111110100111110010101111010011",
    592 => "11100011011110111100000100110000",
    593 => "10001111111011110001100010100101",
    594 => "11101110110011110000111110011101",
    595 => "11111101101011110110001010010001",
    596 => "01111110111111110101011101010100",
    597 => "01110111001011010011111010011100",
    598 => "10010011111110010100001011010000",
    599 => "01101101101100010101010100111010",
    600 => "01111110111111111001111011010111",
    601 => "11111111010000111001110010011000",
    602 => "11000110111111111100100111111100",
    603 => "10001111111011000111110001010100",
    604 => "10110101111110010110101001001100",
    605 => "01111001111111110001010000101111",
    606 => "11111101101111110101111010011001",
    607 => "10111111111111111110110101111101",
    608 => "01110101111111111110110111000111",
    609 => "11111110111101101100100100111000",
    610 => "01101110011011111001000110101000",
    611 => "01101111111111101011110111100000",
    612 => "11101111101111110001010100010000",
    613 => "11110100001111110011011011101010",
    614 => "11100101111111111000110000010010",
    615 => "10111000010000111010000010011010",
    616 => "01101011011111110101101100101001",
    617 => "01001110111011011111101101111000",
    618 => "01100110111111100000100110100111",
    619 => "01100111001101110111010101010110",
    620 => "01111110111111111011111000111000",
    621 => "10110100011111010011010100111110",
    622 => "01101110011010110000101100101101",
    623 => "11111110011111110011010001001100",
    624 => "10111111011111110110110100001111",
    625 => "11111011101010111010011000011010",
    626 => "01001111101111101000110001111110",
    627 => "11101111101111111001100101100100",
    628 => "11111010011001100110100100010011",
    629 => "01101110110111111010000101101001",
    630 => "11111100011010111011010011100110",
    631 => "10111110111011010110110100101010",
    632 => "11101011010111110011110100011111",
    633 => "10110110011101111111011111100000",
    634 => "11110110010110101011001000011101",
    635 => "11101111101111010011001000110001",
    636 => "01111111010111101010010101110111",
    637 => "11100111111011111101011111011000",
    638 => "01111101111100101000010100000011",
    639 => "01011011111101011100000100001100",
    640 => "01011110011110101100010010100110",
    641 => "11011111110101110000101011010110",
    642 => "10111111101111011001001001000100",
    643 => "11011100101100100111111001001010",
    644 => "01111111011010111010101001110111",
    645 => "01011111110111001000001010000101",
    646 => "01111111011111110111110111010111",
    647 => "11101101100111001001101111010010",
    648 => "01111011111010101111110100010010",
    649 => "10010110000101010100110101101110",
    650 => "01011111011110111111000110011100",
    651 => "11110111110011101001001110010110",
    652 => "11111101101111100110100011101010",
    653 => "01110111110111011110001111111011",
    654 => "01111111010001010010011101001111",
    655 => "10111111110100110011001101111110",
    656 => "11111001110011100111010110101111",
    657 => "01110000001011111000101001010001",
    658 => "01011111110111110010011111110011",
    659 => "01010110011111100111110010111010",
    660 => "11111011110100110100100011001111",
    661 => "01111011011110111011001010101010",
    662 => "01001111111111100001110111100000",
    663 => "01111011111111111111100011111110",
    664 => "01011111011111001100001000100111",
    665 => "01111000111111110101010011100111",
    666 => "10111101110101110110101000000110",
    667 => "01001111100110011011110101011101",
    668 => "11100110101011010011000110010010",
    669 => "01100101001101001100010001000001",
    670 => "01111011111101111001111011101101",
    671 => "01111001111111110001011011011001",
    672 => "00111111110011110101101000010110",
    673 => "11011110110101110011011000010110",
    674 => "01001111101111111101000101100010",
    675 => "11111111011111101111001001011111",
    676 => "11111011010111011001010000101000",
    677 => "01111111011011110000101000110101",
    678 => "11110111011111110011000111001001",
    679 => "11111110111110100000101000010011",
    680 => "01111111010110111101011111011011",
    681 => "10011111111111010100010010000010",
    682 => "01110111111101101100001000011010",
    683 => "11101111110111110111100111100101",
    684 => "11110011111111101100000001001100",
    685 => "01111100111101110011000011001010",
    686 => "11101111111011011111000100110100",
    687 => "11111011100101101111011100001101",
    688 => "11111111011111010000100101111000",
    689 => "11011101101111111011000111011001",
    690 => "10111111110111101101010011001001",
    691 => "01010111101110101111001111110000",
    692 => "11111110010000110110001101001011",
    693 => "01111011011011101000110101000011",
    694 => "11110111111001110111001000011100",
    695 => "01110110101101111101000001011111",
    696 => "01101011011101000100011111011001",
    697 => "01111110110111110110001100010110",
    698 => "10110101001110000001010011111100",
    699 => "01000101110111111001010101000010",
    700 => "11001111011101100001110101001111",
    701 => "11111011111111111111110111001000",
    702 => "11011010100110111011000010101011",
    703 => "10100110110110111011011011110011",
    704 => "01111010001111101101100100100100",
    705 => "01111110011111111010001010011110",
    706 => "11100001000011110100100011110000",
    707 => "11011011011111111010001100000100",
    708 => "10111011011111110111111001100010",
    709 => "01011011111101010111100001000110",
    710 => "10011111111111111111110111000111",
    711 => "11100011011001101010100111110010",
    712 => "10100111101111110001101001100100",
    713 => "11101111010011111101111000001100",
    714 => "10111111111111110111101001001100",
    715 => "01111011111110010110111110101010",
    716 => "01110111010110001010111100111110",
    717 => "01011100101100111011100111010111",
    718 => "11111011111001110010011100000010",
    719 => "01101111111110110010101001100111",
    720 => "11110111111111110110110110001101",
    721 => "11101101111101011100110100001101",
    722 => "11001010111101110000010101111011",
    723 => "10111111110101010111101101101010",
    724 => "01100111111001001011011110100001",
    725 => "01110111110010111111010111000111",
    726 => "10100111000001111001101011010100",
    727 => "01110111101111110011100110010011",
    728 => "01100110110101111010100110101000",
    729 => "11011101111111110100011010101111",
    730 => "10111000101110001101000010000111",
    731 => "01111011111111010110111001111110",
    732 => "11111100100111001100110111000101",
    733 => "11011010110111110011010111010100",
    734 => "00111111111100101100000111100000",
    735 => "01011111111111110110001010100110",
    736 => "01101111101111110010010001100111",
    737 => "11011111010010011011111001101001",
    738 => "11111101001101110111011100100010",
    739 => "00111111111101100101100100110110",
    740 => "10101111010110111001110101111011",
    741 => "01101110110010111101011011101110",
    742 => "01100111011011010110011000001010",
    743 => "11110111110101000010000101111001",
    744 => "11111111010110011100111010100011",
    745 => "01111111011010110010001100100100",
    746 => "11111110101010110010000010100011",
    747 => "11101111111011010110110000100000",
    748 => "11110110100001110101101110101011",
    749 => "01101111001010110110110010010000",
    750 => "01101111111000111100111001000110",
    751 => "10101110111011101010110011001010",
    752 => "01101110110011110010101001011011",
    753 => "10111110001111111011100001001000",
    754 => "01101111011010010100011010110111",
    755 => "01111000011100001110100111101111",
    756 => "11111010101100110101001000011101",
    757 => "01111111010101010100101110001001",
    758 => "01111110111011101110110011011100",
    759 => "01111010111111010111001101001011",
    760 => "10101011011111011110100110000100",
    761 => "01110111111000011101111011001110",
    762 => "01001011001111101010101110001001",
    763 => "01110101010011110000101001110100",
    764 => "01011101001110111011000110111100",
    765 => "11111011101010111101111110011000",
    766 => "00111111111101111011100101011011",
    767 => "01001101101110111010011011110110",
    768 => "01111001111011111001101000010110",
    769 => "11100111111110101110100100111001",
    770 => "11111010110101110000001100000010",
    771 => "11011111111111011101100110101110",
    772 => "11011111111011111000100110010111",
    773 => "01101000011101111101100001101111",
    774 => "10000011111110110001001001100111",
    775 => "01111100001111110111111110010110",
    776 => "10011110110110111100110011111110",
    777 => "01100001101110110101011000001011",
    778 => "11111101011111010110001001010101",
    779 => "11111100111011110001011101000011",
    780 => "01110001101011011000000000000110",
    781 => "01111011101111011101001011000001",
    782 => "01011100111111010010111110101110",
    783 => "01001001000111101111100101011011",
    784 => "01111110110111011000110000010110",
    785 => "01011111111111111011001001010001",
    786 => "01111111011111110011110011111111",
    787 => "01111101111111010100010001000101",
    788 => "10011011110101110000011000001001",
    789 => "11111011111101100010101100111000",
    790 => "11001111100011101001011101010001",
    791 => "10101111101101011000110111110100",
    792 => "11101010111111111000100111111010",
    793 => "10001111111100110100101011111100",
    794 => "01111110111011110110001110110101",
    795 => "01111101101111001101111000101011",
    796 => "11101111111110011000001011001001",
    797 => "01110111111011001101100100110111",
    798 => "01010111111110110110001111110011",
    799 => "10111100011111000000101100000111",
    800 => "11001101111011010100001010001000",
    801 => "11011011110111011010001010000111",
    802 => "10100100010110011000100001101110",
    803 => "01110111111111000001101101110010",
    804 => "01111110111111111010111001001001",
    805 => "01110101111111111011100101010011",
    806 => "11011111111111111110000100011001",
    807 => "01101111111110110110111100001111",
    808 => "11110111111011110011101001101000",
    809 => "01011111101111110111001011000010",
    810 => "10001111110011100001101111100110",
    811 => "11111010101011111110010011011001",
    812 => "01000111011101110010100000010001",
    813 => "01111010100110011011101100111111",
    814 => "01011101110001101101001100100001",
    815 => "11111111011111100100010001110010",
    816 => "11001100111110111000111001000001",
    817 => "01100100011101110000010001100001",
    818 => "11111101101101100001000000100001",
    819 => "11110001001111110101001000000000",
    820 => "11110001011011110101010100110010",
    821 => "11011111111111100101010100011101",
    822 => "11101111110111111001100011110001",
    823 => "10110100111111111010001100111001",
    824 => "01111111011111000101010100101101",
    825 => "01111100110101111110110010001111",
    826 => "11101111110011111000000001100111",
    827 => "01011011101111011100011101011010",
    828 => "00111111111011010000010110010100",
    829 => "10011011110111110100000011111001",
    830 => "11011011101100111101100010101101",
    831 => "11011101000111100011110110001000",
    832 => "01001111111010010001001010110011",
    833 => "01100110101110111001101011000010",
    834 => "11101111111101110011111011100100",
    835 => "10011111111101110010010111000010",
    836 => "11111011101011110111001110001010",
    837 => "01111001111110011110101100010101",
    838 => "01111011011111010000010011111011",
    839 => "11011110110111011111100110000110",
    840 => "11111111010111111011111100000110",
    841 => "10110111110111111001001011101111",
    842 => "11010101111101111101001010110000",
    843 => "11111111011110111000110111011101",
    844 => "01101000111000000001111000100001",
    845 => "01111101101001110100101000010110",
    846 => "11011011001101101111000100000111",
    847 => "01011100111011010010111010001011",
    848 => "10101011100101011011101011101101",
    849 => "11101011000011010100101001001111",
    850 => "01001111111010110111000111001111",
    851 => "11111011111001110110101001110000",
    852 => "11101110010101011010010010010000",
    853 => "01111011111000100100100011111110",
    854 => "10110100010111100000101111000111",
    855 => "10011110111011100101011000110011",
    856 => "11100011111100111110011011001011",
    857 => "01111000101110110110110111110100",
    858 => "11010110111111101110111111001101",
    859 => "01111110011101011101011000001111",
    860 => "11111101110111101111111100101110",
    861 => "10110011111111110010101111000001",
    862 => "11111001100111111100111111011110",
    863 => "11011111111000101101011000101011",
    864 => "01111011001110111110010110010001",
    865 => "01101111111011111011000100111100",
    866 => "01110110110111101010010011011011",
    867 => "11111100101000100110100010010101",
    868 => "01010101001000110111011101010111",
    869 => "01011111111101110111010001101010",
    870 => "11111010010111111110000110100011",
    871 => "11111011111100001011011010111101",
    872 => "01111011101011111010010011011100",
    873 => "11011101100110111010100100010000",
    874 => "01011101111111111100111001101010",
    875 => "11111011111111011100111111101010",
    876 => "11011111011101111000011100101110",
    877 => "01111101101010111110001010001011",
    878 => "01001011001011001011011111110101",
    879 => "11110110111111011101110010101100",
    880 => "01010101110101110011101010100100",
    881 => "11111111001111101110010000000001",
    882 => "11100101111101001011001000100101",
    883 => "01101101111011111001000101101100",
    884 => "11011100111011011011000100110100",
    885 => "11001111110011110110000101110011",
    886 => "01101111110111010100101000100110",
    887 => "00111111110101010010010110111100",
    888 => "10101111111010111110001111011001",
    889 => "01111011101011011101100011110100",
    890 => "10111111101101000001000110000101",
    891 => "01101101101010111111011000001110",
    892 => "11111011100111110000100110100011",
    893 => "11111110111101111001111110110100",
    894 => "00111111110110010010010010101011",
    895 => "01111100111110001010101010111011",
    896 => "11111010101111111001010011011110",
    897 => "11110111111101011000100111011110",
    898 => "11010111010111001100101010000001",
    899 => "11111110011111010010011000101111",
    900 => "01001010101111001110111000010101",
    901 => "11001101011111011001110100101000",
    902 => "01111111011111111101000001101101",
    903 => "11111101111100111101110001111001",
    904 => "11011011101111110010101110111100",
    905 => "01101101111101111010110010010111",
    906 => "01001110011011111111000100100111",
    907 => "01111000111110111000001100010100",
    908 => "01111101110011110001111000010000",
    909 => "10111111111111101110110100000011",
    910 => "01111110111111110010100010001001",
    911 => "11111011000110111010100101000000",
    912 => "11101111111111110100101011100110",
    913 => "10101101011011111101100101110111",
    914 => "11101111111011111100001001001000",
    915 => "10011111111001101111011010001011",
    916 => "01111101111000000101011110100110",
    917 => "01001001110111111110001101001000",
    918 => "10011011010100010110101000101011",
    919 => "11111111001111110101111010100001",
    920 => "01111110111110010001001000100011",
    921 => "01110011100110110010111110011111",
    922 => "11111011111111110111011000001000",
    923 => "11101100111111100011011010100010",
    924 => "10001011111001111111100111101010",
    925 => "10111100111111101001101001011001",
    926 => "11011000111101110010101110101011",
    927 => "10110111101100110101101011110100",
    928 => "11011101111111111011001100101100",
    929 => "01010111110011001110101000011110",
    930 => "01110100010010100101001110100000",
    931 => "10110110110001111110111000000000",
    932 => "01011101100111000010111011110010",
    933 => "01111110101110101111111101001010",
    934 => "01110101010101111010000000110000",
    935 => "11011110111111100011011101110001",
    936 => "11011111111011010011011001000001",
    937 => "11001011111101110110000110000110",
    938 => "10001111011111111110110001011110",
    939 => "01011111110100110001101111111001",
    940 => "11011111111011110100010010110100",
    941 => "11110110111111110001001110010000",
    942 => "11111101101111111101100111111000",
    943 => "11111000111010110101000111111001",
    944 => "10010011111111101101111111011010",
    945 => "01011110111111111111100100001111",
    946 => "11111010011110111111000000011011",
    947 => "11111001010110110110110101011110",
    948 => "10101110110100000110110110101100",
    949 => "11101011111111110110011100011110",
    950 => "11100110001111101101010000011001",
    951 => "11110110011111111110001011101111",
    952 => "01111111011110111100111000001110",
    953 => "11111110111001100110111000100110",
    954 => "01111011001101100001100100001001",
    955 => "01101111110101111101010110011110",
    956 => "10110111011110000111000111111101",
    957 => "01111011011011101111111010000101",
    958 => "01111011101000110110001101100110",
    959 => "11011011000111110111111011101011",
    960 => "11111110001011011101011001110011",
    961 => "01001011000110110011110111100011",
    962 => "10111100011010110000100110010001",
    963 => "01010001011111110001111110111011",
    964 => "11101111110011010110110001011011",
    965 => "11111010100110100010110010110110",
    966 => "01110111101111111001010111001111",
    967 => "01111111011111110101001110010100",
    968 => "11100101101100111011000011000010",
    969 => "11111111011001110010000011100110",
    970 => "11110101101011110011000010011110",
    971 => "10010110101101001001110111100111",
    972 => "00111111110111110001011011001110",
    973 => "11011110011111110000001011011100",
    974 => "01100100111111110100100001000101",
    975 => "10011101010111110010001100110001",
    976 => "10111101110011010011110110111111",
    977 => "11101011100110110011111000011110",
    978 => "01101010111101010110111100010110",
    979 => "11011011111110011011000010010011",
    980 => "01110101111101110111000001010010",
    981 => "10110111111111001001110111000010",
    982 => "11101110111111100001000010011100",
    983 => "10111111101110110111011001100011",
    984 => "10101111001101100110001001100100",
    985 => "11100111011111111100101101010110",
    986 => "11101110001110110111101001110100",
    987 => "11000111101111011010000110010010",
    988 => "11011100110010110000111011110001",
    989 => "01110101100001110100110000011000",
    990 => "10111001111110111111000110000101",
    991 => "01101111111011111111000111010000",
    992 => "01111000111111110011001111110011",
    993 => "11111011111110001001101001110111",
    994 => "01011111011011110110010111001011",
    995 => "11111110101111101001000011000001",
    996 => "01101110110111111010110001100000",
    997 => "11111101111111010110011101010110",
    998 => "11011101111110101111110011100100",
    999 => "11111111011001000010011011000011");

  constant ans_lut : lut := (
    0 => "11111011101111011110001101010010",
    1 => "01110111111011111000000000001111",
    2 => "01111011110111100101111001000011",
    3 => "11011101100111011001011110100100",
    4 => "11111101001101111110101111101000",
    5 => "01111111011101101101100000001101",
    6 => "11000000000000000000000000000000",
    7 => "01101111011110101010111110111111",
    8 => "01011110110101100101110010001011",
    9 => "11011010011111101011100010010100",
    10 => "11010011011111101111010011111111",
    11 => "11110111010111001100010101001010",
    12 => "10111111100000000000000000000000",
    13 => "11111100111110111000001001110001",
    14 => "11011110101110111001101011101111",
    15 => "01111111010111011111101001001011",
    16 => "01111011010111111001100111100110",
    17 => "11111011101010101111000100101100",
    18 => "10111111100000000000000000000000",
    19 => "10111111100000000000000000000000",
    20 => "10111111100000000000000000000000",
    21 => "11011110111110110111110100011111",
    22 => "11111011111011110010010101101000",
    23 => "11101110111100101111100011010110",
    24 => "01101111110101011101000000010110",
    25 => "01110110111110111010000100100011",
    26 => "01111111000111110010001111111111",
    27 => "01111110111111111111000100110001",
    28 => "11101111011111111011101001010100",
    29 => "11000000000000000000000000000000",
    30 => "01010011111101010011010001010000",
    31 => "10111111100000000000000000000000",
    32 => "11110000111110001111110010110101",
    33 => "01110111101011001101001111111101",
    34 => "01010001010111111000010110101111",
    35 => "10111111100000000000000000000000",
    36 => "11111011100111101000011011010000",
    37 => "01110110111111101101011000111000",
    38 => "01101011001011111010010011011010",
    39 => "10111111100000000000000000000000",
    40 => "01101101110011100010100101110101",
    41 => "11011010000111110010000100100010",
    42 => "11100100111001000001100101000010",
    43 => "01011101111101110000110111101010",
    44 => "11111010111110111111100001011001",
    45 => "11111101011111100000011011001001",
    46 => "11111010111111111101100100110100",
    47 => "11111111010101010010101111100011",
    48 => "11110011111101011110100001011000",
    49 => "10111111100000000000000000000000",
    50 => "01011011101111111011110011100110",
    51 => "01101111111010110010011101101100",
    52 => "11011011110110110010010010101111",
    53 => "01001110111101001111011111001011",
    54 => "01101001111100110001000000111111",
    55 => "10111111100000000000000000000000",
    56 => "10111111100000000000000000000000",
    57 => "11110111101110111010101010111001",
    58 => "11111110111011001001000100000010",
    59 => "11111110111001110100111100001100",
    60 => "10111111100000000000000000000000",
    61 => "10111111100000000000000000000000",
    62 => "01011111111111110100101100100110",
    63 => "01111010100100111011101101111001",
    64 => "11111000011111111100000010011110",
    65 => "10111111100000000000000000000000",
    66 => "11000000000000000000000000000000",
    67 => "11000000000000000000000000000000",
    68 => "11100111110111100101110010110101",
    69 => "01110011111010100100010001010011",
    70 => "11111110111111000110001111010011",
    71 => "10111111100000000000000000000000",
    72 => "11110011011101011010101110000010",
    73 => "11011100111111100001111001001011",
    74 => "01111001011100011011110100010001",
    75 => "01111101101111101110101100011010",
    76 => "10111111100000000000000000000000",
    77 => "01111111011101010101100010110011",
    78 => "10111111100000000000000000000000",
    79 => "01110111111111011011111101111100",
    80 => "10111111100000000000000000000000",
    81 => "01110010110001001100010000100010",
    82 => "01011011011101010101111011000101",
    83 => "10111111100000000000000000000000",
    84 => "11111011111111111111011110000001",
    85 => "11111011111110011010101011111011",
    86 => "01011110011111101010110010011100",
    87 => "11000000000000000000000000000000",
    88 => "01111010111110110111000110011010",
    89 => "00111111100000000000000000000000",
    90 => "11100110111111101010011100110110",
    91 => "01011111100101011100100111011111",
    92 => "11101101010110111000011011101000",
    93 => "01101100011111110101001110001011",
    94 => "11000000000000000000000000000000",
    95 => "01011111101010110101101111100110",
    96 => "01000110111111011111111000000000",
    97 => "11111110111101111101000100011100",
    98 => "01001111110010110101110101011111",
    99 => "11111110111111110100000111010110",
    100 => "10111111100000000000000000000000",
    101 => "10111111100000000000000000000000",
    102 => "01101111101111010100101100101000",
    103 => "10111111100000000000000000000000",
    104 => "01111011100110100111100000100000",
    105 => "11100111110111001011011001100000",
    106 => "11010110111010110000000100011111",
    107 => "01111101001001011110101101110001",
    108 => "11111101111011101110111000100101",
    109 => "10111111100000000000000000000000",
    110 => "11010111010111101001010011000010",
    111 => "11110110100111001100110100001011",
    112 => "01110111111011111001000001000000",
    113 => "11011111111111100011101110001010",
    114 => "11101110111100110110001011111110",
    115 => "01110010110111110011001011000001",
    116 => "11110111101111111101101111001000",
    117 => "11101100111011000000001100110011",
    118 => "01111110101000110100101010000101",
    119 => "01101111101111110101001010000101",
    120 => "01000110101110101010100000000000",
    121 => "01011111100101010011011101100101",
    122 => "11111100101101111111111111101011",
    123 => "11011100111111101100110111010111",
    124 => "01111110101110011010001011000000",
    125 => "11011110110010100000001011000110",
    126 => "01101101111001111110101111111110",
    127 => "01011110101111111000110011111011",
    128 => "01111011110000111001011001011110",
    129 => "01011110111111001111011001000101",
    130 => "11111011011110011000111110110011",
    131 => "10111111100000000000000000000000",
    132 => "11010110111101111101000101011001",
    133 => "01101011111111101101110110001010",
    134 => "11001111101101100010010010001100",
    135 => "01111011111110010110010010001000",
    136 => "01111101011111111001001011000101",
    137 => "01100111111111110010100000011001",
    138 => "11111011111110110011000101101010",
    139 => "10111111100000000000000000000000",
    140 => "11000000000000000000000000000000",
    141 => "01101110101101111000111011000111",
    142 => "11111110011010111011100100110000",
    143 => "01101101111111101000001111101100",
    144 => "01010101111011010110100000001110",
    145 => "01010101111111110000010011110000",
    146 => "11101101100011110100001000100000",
    147 => "00111111100000000000000000000000",
    148 => "01000101101111110010100000000000",
    149 => "11110110100010100101011110100001",
    150 => "01011001111011111011000111000010",
    151 => "10111111100000000000000000000000",
    152 => "01111110111111111001100011101111",
    153 => "11011111110111111111111001001010",
    154 => "01110111111111111000010010010110",
    155 => "01110001111111111100011101011011",
    156 => "01011100110111010101010100011011",
    157 => "11010111011111111010111011110101",
    158 => "01111111001101111111101001010000",
    159 => "01111011101100010000101011000101",
    160 => "11111011111111111110110000001001",
    161 => "11101111110101011111010000101101",
    162 => "01101111001011110000011010101011",
    163 => "11111011011111011110001001011000",
    164 => "10111111100000000000000000000000",
    165 => "11101110111001010111110011100010",
    166 => "01001011111111010101101000101101",
    167 => "01100011111010110010011000101111",
    168 => "01111001101100110001001010000101",
    169 => "01011111010010100110111011110101",
    170 => "01011010111111111101101101010011",
    171 => "01101111110111111100111111001001",
    172 => "11010111111101110110111110100000",
    173 => "01110110010110110101101101011100",
    174 => "10111111100000000000000000000000",
    175 => "01010110111101110100010100100110",
    176 => "01111011111111110000111001100110",
    177 => "01101010101111111010010001011101",
    178 => "11101011101111010100110101010111",
    179 => "10111111100000000000000000000000",
    180 => "11111011111111110100010111010111",
    181 => "01111110010111011010000000000011",
    182 => "01111101111001010111010110100111",
    183 => "01001101011110110110100111110111",
    184 => "11011111100111111010101111101100",
    185 => "01110111101011110100111111100010",
    186 => "01111110100111110100010011111101",
    187 => "11101110011111111100010010100100",
    188 => "10111111100000000000000000000000",
    189 => "11111111001110010111111110111111",
    190 => "01111110110110010100011110101011",
    191 => "11010001110110101110111010101010",
    192 => "01111111010011111100101000110111",
    193 => "01101011111010111000110011011110",
    194 => "11110110111111100110011110101110",
    195 => "01110011100110110100011111110111",
    196 => "01111111010111101011111010010110",
    197 => "01111111011110010001101011100011",
    198 => "01001011101011101000110100010011",
    199 => "11101111100011001000110111100000",
    200 => "01111100100011101110100110001011",
    201 => "11000000000000000000000000000000",
    202 => "10111111100000000000000000000000",
    203 => "10111111100000000000000000000000",
    204 => "10111111100000000000000000000000",
    205 => "01001011010000011100011100011010",
    206 => "11101001111111111101100111000101",
    207 => "11111011110011110100000111011110",
    208 => "01101011111001111010100000111110",
    209 => "11010101011011100011100110010001",
    210 => "01111011110011010100001000100000",
    211 => "01101011111010111111101011110110",
    212 => "01010111111111111010000000001110",
    213 => "01010001011110111110000101000010",
    214 => "11011111111101101001111110010011",
    215 => "01110111111000000110000101111110",
    216 => "11110010101101110001101000110101",
    217 => "01111101010110111001000001010000",
    218 => "11110101100101101000011111110101",
    219 => "01011101111110011011110111111100",
    220 => "11100111101011110010101111001000",
    221 => "01111101101010101000100000111111",
    222 => "11111010000111100011001001000110",
    223 => "11110001111110100000111111110001",
    224 => "10111111100000000000000000000000",
    225 => "01111101111111111001000010111110",
    226 => "11101110110111111101000011000010",
    227 => "01110111010110010110000100000011",
    228 => "01111011111111100001101000111010",
    229 => "10111111100000000000000000000000",
    230 => "01111110011110101101011101001100",
    231 => "01011111011010111110001100011000",
    232 => "10111111100000000000000000000000",
    233 => "01111000110111100111110011011010",
    234 => "11000000000000000000000000000000",
    235 => "11001111111111101010011100001000",
    236 => "01101111011010111001111100100101",
    237 => "11111011111110111101101000000100",
    238 => "11111011111111100010100101010110",
    239 => "11110001110100111001001010110110",
    240 => "01101111111101111001100101111010",
    241 => "01101111001111110000100111001110",
    242 => "01101011111111010000110000001110",
    243 => "01111110111100111110011000001001",
    244 => "11111101010101011101000011010010",
    245 => "10111111100000000000000000000000",
    246 => "01111011111111110001110010010110",
    247 => "11011111011101110101010011111110",
    248 => "11111110011110011001000110001011",
    249 => "11111110111011101100001100101010",
    250 => "11111111001011110110011111011100",
    251 => "10111111100000000000000000000000",
    252 => "01011010111111001000011100100100",
    253 => "01110111101111110111001000110101",
    254 => "01111100101011110111111000100100",
    255 => "10111111100000000000000000000000",
    256 => "11011101111111111011000001111010",
    257 => "11101101010111001010011001001011",
    258 => "10111111100000000000000000000000",
    259 => "11101111110011010011010100110110",
    260 => "10111111100000000000000000000000",
    261 => "01111110111100010100000000111010",
    262 => "11010111111001011000000001100101",
    263 => "01000111110111110111111100000000",
    264 => "11110111001111111000111000110010",
    265 => "01010111011011111110000010111101",
    266 => "01110111111111110111100001100010",
    267 => "11101110100111111011000011011100",
    268 => "01111111001101011000100010000001",
    269 => "01110011110111110110011010011010",
    270 => "01111101111111101011100100110011",
    271 => "01111101101011110011101010110100",
    272 => "11111001001001110001101001001011",
    273 => "11111101111111101110101011111010",
    274 => "01111101111111010100101101001000",
    275 => "10111111100000000000000000000000",
    276 => "11110101110110010010001100100110",
    277 => "01111111001101111101011100110001",
    278 => "11111100111111111011011011111001",
    279 => "11111101110011111110011101100011",
    280 => "11101101111101110101001011010111",
    281 => "10111111100000000000000000000000",
    282 => "01011010111111100000101001000100",
    283 => "11110101001111110110111010001011",
    284 => "11111111011011111010110011111100",
    285 => "11111000011011100001010101110000",
    286 => "11000000000000000000000000000000",
    287 => "11110111111111111110101010100001",
    288 => "01111110111111110110110111100001",
    289 => "01000111110111110101100000000000",
    290 => "01011111111011011010100000010010",
    291 => "11011110111100000001100000101110",
    292 => "11111111011111010110111110010101",
    293 => "01011101111001111010000000100111",
    294 => "11000000000000000000000000000000",
    295 => "11101101111111010110011001000101",
    296 => "11011101111010110000101110000110",
    297 => "11101111011111010111010011110001",
    298 => "01011111100111100101101111001010",
    299 => "11011011111111110011011000111011",
    300 => "11000000000000000000000000000000",
    301 => "01111110110111110000111010111110",
    302 => "10111111100000000000000000000000",
    303 => "01101110111110111011111110101011",
    304 => "01011110101110110111001000110100",
    305 => "11101101111110110000011000001100",
    306 => "11100110011111000100111110001111",
    307 => "11111110111111010011111110010001",
    308 => "11000000000000000000000000000000",
    309 => "11111000111010111011101111101101",
    310 => "11010101100111111010010101100110",
    311 => "11111110110110110101001111101100",
    312 => "10111111100000000000000000000000",
    313 => "10111111100000000000000000000000",
    314 => "01110110111101101001001100010101",
    315 => "01111011111100010100001000101001",
    316 => "10111111100000000000000000000000",
    317 => "11010111101110011011100110110010",
    318 => "11111010111110110111101110001110",
    319 => "11110100010011110001011110001110",
    320 => "10111111100000000000000000000000",
    321 => "01011101111111101011101001011010",
    322 => "11111110100101110110011010111001",
    323 => "11111001111011110111011101000110",
    324 => "10111111100000000000000000000000",
    325 => "01110100111110110100110010010000",
    326 => "11111001101111101111111000000101",
    327 => "11011101101011111101100110101100",
    328 => "01110111011111101101101111101111",
    329 => "11110111100011000101011111101000",
    330 => "01101111011111101000100111100001",
    331 => "11010111011101110111011010010000",
    332 => "10111111100000000000000000000000",
    333 => "11011011111101110001001010010001",
    334 => "11001101110111001001011110110111",
    335 => "11101110101111101100010110110110",
    336 => "11111111000101111001001100011100",
    337 => "11111111011001110000111111001001",
    338 => "11001111101101110111110010100010",
    339 => "01101111111111110010111100011110",
    340 => "11000000000000000000000000000000",
    341 => "11111011110111111111000011111000",
    342 => "11001111111110101101011010011000",
    343 => "01111011110011101100110111010100",
    344 => "11110011011011110110100100000110",
    345 => "11111101111111000110101000111101",
    346 => "10111111100000000000000000000000",
    347 => "01110010111011111101111110101011",
    348 => "11111111011111100101111010011001",
    349 => "01001011111110111111110101000011",
    350 => "11011001001110111010001001010110",
    351 => "10111111100000000000000000000000",
    352 => "11111011111001110000101011001011",
    353 => "11111101111110011111010000010110",
    354 => "11111101100011100111011110001111",
    355 => "01001110101111010100000010111101",
    356 => "01001111111001111000100111101110",
    357 => "10111111100000000000000000000000",
    358 => "01111111001101010001000000100011",
    359 => "11011111110111000101111100000001",
    360 => "01111110111011110000011010111001",
    361 => "01100101111110111100001000011010",
    362 => "11011111101111110010111000100000",
    363 => "01111111011011110111100011110101",
    364 => "01011111011010111101100111011011",
    365 => "01111100101111110000001101110111",
    366 => "11010111111111110100111010000000",
    367 => "11101111011110001011101100111011",
    368 => "01110011000101010001010000111000",
    369 => "11111110011101100000101010001010",
    370 => "11111011110100110011000001111011",
    371 => "11011110111001000101001010110110",
    372 => "10111111100000000000000000000000",
    373 => "01001011111111010010011011110100",
    374 => "01101011011110110101001100000011",
    375 => "11111110111101011000100001101100",
    376 => "11111110111111110011100010101101",
    377 => "11110011111011111000101000111011",
    378 => "01101100111111001001110011111101",
    379 => "10111111100000000000000000000000",
    380 => "11111111011011010010011000000101",
    381 => "01011110100010000100111101011011",
    382 => "01100111111111001001011100011110",
    383 => "01110111111011010000110111100010",
    384 => "11011011011100111010000000010011",
    385 => "01011110111101100001100110010101",
    386 => "01011011110011111101011011100011",
    387 => "01100000111110101101111000100100",
    388 => "01101100111111111011011010101110",
    389 => "01111011111011110101010011011001",
    390 => "01001111101111110110110101001111",
    391 => "11000000000000000000000000000000",
    392 => "01011100111110110011111100101000",
    393 => "11101010111100101101001101011010",
    394 => "11110011011111110111100110111010",
    395 => "01011011111011011111100000111111",
    396 => "01010011110111101011110010001111",
    397 => "10111111100000000000000000000000",
    398 => "10111111100000000000000000000000",
    399 => "11111011110111011111100011000001",
    400 => "11110110111101111001010001110000",
    401 => "01001111001111110001101001111101",
    402 => "01101111110111100011111101000101",
    403 => "11101100110111011001111011001001",
    404 => "10111111100000000000000000000000",
    405 => "11110011011110100011111111101001",
    406 => "11001011101111110010011001010000",
    407 => "10111111100000000000000000000000",
    408 => "10111111100000000000000000000000",
    409 => "01111011100011111011100111010111",
    410 => "01111011011110111011010011000011",
    411 => "01111010011111111111110001111100",
    412 => "11001111111001110100000110101100",
    413 => "01011011001111110100011101010010",
    414 => "01110001111111110001000101010011",
    415 => "01111011100111011010011001011101",
    416 => "01100111101111101101000100100110",
    417 => "10111111100000000000000000000000",
    418 => "00111111100000000000000000000000",
    419 => "11111000111111110111100001110010",
    420 => "10111111100000000000000000000000",
    421 => "01010011100101111010101111110100",
    422 => "01111001111111110011111011001100",
    423 => "11111110111101111011010001110101",
    424 => "01111011111111111100000101111010",
    425 => "11111101111101100010101100011110",
    426 => "01111101110010100111101101010111",
    427 => "01001010001001110100101110111100",
    428 => "11010011110111111010011100111000",
    429 => "10111111100000000000000000000000",
    430 => "01111011110110011111010011011110",
    431 => "11010111101001110000100100100100",
    432 => "01111011111111110100101100111100",
    433 => "11010011111011110100001101101010",
    434 => "11111011001111110101001001101100",
    435 => "10111111100000000000000000000000",
    436 => "01111000001111110101011011010000",
    437 => "01011111011111101001100111100000",
    438 => "11111100111111101101100101110100",
    439 => "01111100110010111101011001000000",
    440 => "11111101011000111001011011110001",
    441 => "01111101111111111011010100001100",
    442 => "11101001111110111001000110001100",
    443 => "10111111100000000000000000000000",
    444 => "01100111111111110110111111101111",
    445 => "11000000000000000000000000000000",
    446 => "11111100011111010111001010110101",
    447 => "11110111111010110111111011011010",
    448 => "11100001011110111000111010101101",
    449 => "01001010011100111100001110000000",
    450 => "11011111101000110011001010011100",
    451 => "01111101111111011011010000110011",
    452 => "01111111010011011000100111010000",
    453 => "11111101101111110001100001101101",
    454 => "11000000000000000000000000000000",
    455 => "01101011110111110001010100001111",
    456 => "11010111110101110111011011111101",
    457 => "01110111110011011011001111111101",
    458 => "10111111100000000000000000000000",
    459 => "10111111100000000000000000000000",
    460 => "10111111100000000000000000000000",
    461 => "10111111100000000000000000000000",
    462 => "11110010110111101000100100101000",
    463 => "01110110111110110001001001111100",
    464 => "11101101111001101110010001011010",
    465 => "10111111100000000000000000000000",
    466 => "01010101011101111111010101100110",
    467 => "01011110011111011010111011000011",
    468 => "01101101111010010110101000010001",
    469 => "01110110000110110101011101101011",
    470 => "10111111100000000000000000000000",
    471 => "11011111111111111100101111110001",
    472 => "11111110101111010100101000111100",
    473 => "11110011011011000010100010111100",
    474 => "00111111100000000000000000000000",
    475 => "11111111011111111110011001011101",
    476 => "11110011100111110110011000100010",
    477 => "01111010111111010010100011000001",
    478 => "11000000000000000000000000000000",
    479 => "01111111011111110100011010001001",
    480 => "10111111100000000000000000000000",
    481 => "01010110100111111010000100111000",
    482 => "11111001101110110101110110011101",
    483 => "11110011101111011010110010100110",
    484 => "10111111100000000000000000000000",
    485 => "11100111110011010010000100100101",
    486 => "01101011011111110010110000001101",
    487 => "01010100110011111101110001010110",
    488 => "11000000000000000000000000000000",
    489 => "01110101001100111001000000000011",
    490 => "11111111011111011010011000010000",
    491 => "11101110111111110001100000110111",
    492 => "11101110111111100100000010100010",
    493 => "01001101111111111101001111101000",
    494 => "01011011111110110111011100001011",
    495 => "01111011101111111000100011001110",
    496 => "01111111001011111100101100001011",
    497 => "11111011111111101100011011110011",
    498 => "11111011100000110001101001010010",
    499 => "11110110111110100011010101011100",
    500 => "01111110011001110100011111001011",
    501 => "11110111110111111011000001010001",
    502 => "01110111011111101001100101000101",
    503 => "10111111100000000000000000000000",
    504 => "11111101110111110111111001101010",
    505 => "11110111111111010001101111101100",
    506 => "11111110101110110010000100010011",
    507 => "10111111100000000000000000000000",
    508 => "11110111011011110000011101000000",
    509 => "10111111100000000000000000000000",
    510 => "11000000000000000000000000000000",
    511 => "01001101010000010111101000010000",
    512 => "11101111111111001000110000100101",
    513 => "11011111111100000011101011101000",
    514 => "11101111011111100010001110001110",
    515 => "01111101111110010100000110011100",
    516 => "01110111111111110110111001001111",
    517 => "11101100111111111000100001000111",
    518 => "11000000000000000000000000000000",
    519 => "01111011011111111110001000101111",
    520 => "01001011110010110100100011101101",
    521 => "01111011110010010000100100010110",
    522 => "10111111100000000000000000000000",
    523 => "11011110100111110111011101000101",
    524 => "10111111100000000000000000000000",
    525 => "01011111011011110111000111111010",
    526 => "11011111011111110001001101000010",
    527 => "10111111100000000000000000000000",
    528 => "00111111100000000000000000000000",
    529 => "11101111111111110110111001001100",
    530 => "01011000011111111100001111100100",
    531 => "01101011011001110101001110111110",
    532 => "11111011111011110010010001111110",
    533 => "11011111111111110111001100010000",
    534 => "11010111110111110101000101110000",
    535 => "10111111100000000000000000000000",
    536 => "10111111100000000000000000000000",
    537 => "01111111011101111101101011000001",
    538 => "11101110111001001011001010110011",
    539 => "01101011100111010000011001111001",
    540 => "01001100110011010110111110010110",
    541 => "11011111111101110110100111001110",
    542 => "11010110000110110011101010000011",
    543 => "01111111001110110111011010000110",
    544 => "11111111011111111000110010010110",
    545 => "11101101111111110000100100010111",
    546 => "01011010111011110111010001110001",
    547 => "10111111100000000000000000000000",
    548 => "10111111100000000000000000000000",
    549 => "01111111000010111010011110011111",
    550 => "01111111011101110010100100111101",
    551 => "11011011101011001100100101010110",
    552 => "11111011111010011111010100010111",
    553 => "00111111100000000000000000000000",
    554 => "11110110110110010111100001000100",
    555 => "11011111011111110001000101110101",
    556 => "11011101111111111101010000001001",
    557 => "11011111100111111101101111100011",
    558 => "11000000000000000000000000000000",
    559 => "01011001110101101110100000110011",
    560 => "01011111110011110111010001010111",
    561 => "00111111100000000000000000000000",
    562 => "01010011011111101101101111001101",
    563 => "11100101011000110011001100101011",
    564 => "01101110111011111110010100101110",
    565 => "01110111101001110100101110110111",
    566 => "11111101111011111010000100101110",
    567 => "11111011111100100110010001001110",
    568 => "11111110110110110001001101000001",
    569 => "01101111101111111110001001001011",
    570 => "10111111100000000000000000000000",
    571 => "01111011111100011010101010011101",
    572 => "01111000111111010001000110111010",
    573 => "00111111100000000000000000000000",
    574 => "01110111001111111000010011011100",
    575 => "10111111100000000000000000000000",
    576 => "10111111100000000000000000000000",
    577 => "10111111100000000000000000000000",
    578 => "01111101111011010101010101000000",
    579 => "11000000000000000000000000000000",
    580 => "01111111001011011100011111010011",
    581 => "11011001100011011101010000100110",
    582 => "01111110111110011101010100010001",
    583 => "01111001111111010001010000101100",
    584 => "10111111100000000000000000000000",
    585 => "11110101110010110001000111110101",
    586 => "11111011001111110001001011011011",
    587 => "01101011101111110110101111100001",
    588 => "10111111100000000000000000000000",
    589 => "11101111010011110110110000010001",
    590 => "11000101110111100011000000000000",
    591 => "01111110100111110010101111010011",
    592 => "11100011011110111100000100110000",
    593 => "10111111100000000000000000000000",
    594 => "11101110110011110000111110011101",
    595 => "11111101101011110110001010010001",
    596 => "01111110111111110101011101010100",
    597 => "01110111001011010011111010011100",
    598 => "10111111100000000000000000000000",
    599 => "01101101101100010101010100111010",
    600 => "01111110111111111001111011010111",
    601 => "11111111010000111001110010011000",
    602 => "11000110111111111100101000000000",
    603 => "10111111100000000000000000000000",
    604 => "10111111100000000000000000000000",
    605 => "01111001111111110001010000101111",
    606 => "11111101101111110101111010011001",
    607 => "11000000000000000000000000000000",
    608 => "01110101111111111110110111000111",
    609 => "11111110111101101100100100111000",
    610 => "01101110011011111001000110101000",
    611 => "01101111111111101011110111100000",
    612 => "11101111101111110001010100010000",
    613 => "11110100001111110011011011101010",
    614 => "11100101111111111000110000010010",
    615 => "10111111100000000000000000000000",
    616 => "01101011011111110101101100101001",
    617 => "01001110111011011111101101111000",
    618 => "01100110111111100000100110100111",
    619 => "01100111001101110111010101010110",
    620 => "01111110111111111011111000111000",
    621 => "10111111100000000000000000000000",
    622 => "01101110011010110000101100101101",
    623 => "11111110011111110011010001001100",
    624 => "10111111100000000000000000000000",
    625 => "11111011101010111010011000011010",
    626 => "01001111101111101000110001111110",
    627 => "11101111101111111001100101100100",
    628 => "11111010011001100110100100010011",
    629 => "01101110110111111010000101101001",
    630 => "11111100011010111011010011100110",
    631 => "10111111100000000000000000000000",
    632 => "11101011010111110011110100011111",
    633 => "10111111100000000000000000000000",
    634 => "11110110010110101011001000011101",
    635 => "11101111101111010011001000110001",
    636 => "01111111010111101010010101110111",
    637 => "11100111111011111101011111011000",
    638 => "01111101111100101000010100000011",
    639 => "01011011111101011100000100001100",
    640 => "01011110011110101100010010100110",
    641 => "11011111110101110000101011010110",
    642 => "11000000000000000000000000000000",
    643 => "11011100101100100111111001001010",
    644 => "01111111011010111010101001110111",
    645 => "01011111110111001000001010000101",
    646 => "01111111011111110111110111010111",
    647 => "11101101100111001001101111010010",
    648 => "01111011111010101111110100010010",
    649 => "10111111100000000000000000000000",
    650 => "01011111011110111111000110011100",
    651 => "11110111110011101001001110010110",
    652 => "11111101101111100110100011101010",
    653 => "01110111110111011110001111111011",
    654 => "01111111010001010010011101001111",
    655 => "11000000000000000000000000000000",
    656 => "11111001110011100111010110101111",
    657 => "01110000001011111000101001010001",
    658 => "01011111110111110010011111110011",
    659 => "01010110011111100111110010111010",
    660 => "11111011110100110100100011001111",
    661 => "01111011011110111011001010101010",
    662 => "01001111111111100001110111100000",
    663 => "01111011111111111111100011111110",
    664 => "01011111011111001100001000100111",
    665 => "01111000111111110101010011100111",
    666 => "10111111100000000000000000000000",
    667 => "01001111100110011011110101011101",
    668 => "11100110101011010011000110010010",
    669 => "01100101001101001100010001000001",
    670 => "01111011111101111001111011101101",
    671 => "01111001111111110001011011011001",
    672 => "00111111100000000000000000000000",
    673 => "11011110110101110011011000010110",
    674 => "01001111101111111101000101100010",
    675 => "11111111011111101111001001011111",
    676 => "11111011010111011001010000101000",
    677 => "01111111011011110000101000110101",
    678 => "11110111011111110011000111001001",
    679 => "11111110111110100000101000010011",
    680 => "01111111010110111101011111011011",
    681 => "10111111100000000000000000000000",
    682 => "01110111111101101100001000011010",
    683 => "11101111110111110111100111100101",
    684 => "11110011111111101100000001001100",
    685 => "01111100111101110011000011001010",
    686 => "11101111111011011111000100110100",
    687 => "11111011100101101111011100001101",
    688 => "11111111011111010000100101111000",
    689 => "11011101101111111011000111011001",
    690 => "11000000000000000000000000000000",
    691 => "01010111101110101111001111110000",
    692 => "11111110010000110110001101001011",
    693 => "01111011011011101000110101000011",
    694 => "11110111111001110111001000011100",
    695 => "01110110101101111101000001011111",
    696 => "01101011011101000100011111011001",
    697 => "01111110110111110110001100010110",
    698 => "10111111100000000000000000000000",
    699 => "01000101110111111001000000000000",
    700 => "11001111011101100001110101001111",
    701 => "11111011111111111111110111001000",
    702 => "11011010100110111011000010101011",
    703 => "10111111100000000000000000000000",
    704 => "01111010001111101101100100100100",
    705 => "01111110011111111010001010011110",
    706 => "11100001000011110100100011110000",
    707 => "11011011011111111010001100000100",
    708 => "10111111100000000000000000000000",
    709 => "01011011111101010111100001000110",
    710 => "10111111100000000000000000000000",
    711 => "11100011011001101010100111110010",
    712 => "10111111100000000000000000000000",
    713 => "11101111010011111101111000001100",
    714 => "11000000000000000000000000000000",
    715 => "01111011111110010110111110101010",
    716 => "01110111010110001010111100111110",
    717 => "01011100101100111011100111010111",
    718 => "11111011111001110010011100000010",
    719 => "01101111111110110010101001100111",
    720 => "11110111111111110110110110001101",
    721 => "11101101111101011100110100001101",
    722 => "11001010111101110000010101111100",
    723 => "11000000000000000000000000000000",
    724 => "01100111111001001011011110100001",
    725 => "01110111110010111111010111000111",
    726 => "10111111100000000000000000000000",
    727 => "01110111101111110011100110010011",
    728 => "01100110110101111010100110101000",
    729 => "11011101111111110100011010101111",
    730 => "10111111100000000000000000000000",
    731 => "01111011111111010110111001111110",
    732 => "11111100100111001100110111000101",
    733 => "11011010110111110011010111010100",
    734 => "00111111100000000000000000000000",
    735 => "01011111111111110110001010100110",
    736 => "01101111101111110010010001100111",
    737 => "11011111010010011011111001101001",
    738 => "11111101001101110111011100100010",
    739 => "00111111100000000000000000000000",
    740 => "10111111100000000000000000000000",
    741 => "01101110110010111101011011101110",
    742 => "01100111011011010110011000001010",
    743 => "11110111110101000010000101111001",
    744 => "11111111010110011100111010100011",
    745 => "01111111011010110010001100100100",
    746 => "11111110101010110010000010100011",
    747 => "11101111111011010110110000100000",
    748 => "11110110100001110101101110101011",
    749 => "01101111001010110110110010010000",
    750 => "01101111111000111100111001000110",
    751 => "10111111100000000000000000000000",
    752 => "01101110110011110010101001011011",
    753 => "10111111100000000000000000000000",
    754 => "01101111011010010100011010110111",
    755 => "01111000011100001110100111101111",
    756 => "11111010101100110101001000011101",
    757 => "01111111010101010100101110001001",
    758 => "01111110111011101110110011011100",
    759 => "01111010111111010111001101001011",
    760 => "10111111100000000000000000000000",
    761 => "01110111111000011101111011001110",
    762 => "01001011001111101010101110001001",
    763 => "01110101010011110000101001110100",
    764 => "01011101001110111011000110111100",
    765 => "11111011101010111101111110011000",
    766 => "00111111100000000000000000000000",
    767 => "01001101101110111010011011110110",
    768 => "01111001111011111001101000010110",
    769 => "11100111111110101110100100111001",
    770 => "11111010110101110000001100000010",
    771 => "11011111111111011101100110101110",
    772 => "11011111111011111000100110010111",
    773 => "01101000011101111101100001101111",
    774 => "10111111100000000000000000000000",
    775 => "01111100001111110111111110010110",
    776 => "10111111100000000000000000000000",
    777 => "01100001101110110101011000001011",
    778 => "11111101011111010110001001010101",
    779 => "11111100111011110001011101000011",
    780 => "01110001101011011000000000000110",
    781 => "01111011101111011101001011000001",
    782 => "01011100111111010010111110101110",
    783 => "01001001000111101111100101010000",
    784 => "01111110110111011000110000010110",
    785 => "01011111111111111011001001010001",
    786 => "01111111011111110011110011111111",
    787 => "01111101111111010100010001000101",
    788 => "10111111100000000000000000000000",
    789 => "11111011111101100010101100111000",
    790 => "11001111100011101001011101010001",
    791 => "10111111100000000000000000000000",
    792 => "11101010111111111000100111111010",
    793 => "10111111100000000000000000000000",
    794 => "01111110111011110110001110110101",
    795 => "01111101101111001101111000101011",
    796 => "11101111111110011000001011001001",
    797 => "01110111111011001101100100110111",
    798 => "01010111111110110110001111110011",
    799 => "10111111100000000000000000000000",
    800 => "11001101111011010100001010001000",
    801 => "11011011110111011010001010000111",
    802 => "10111111100000000000000000000000",
    803 => "01110111111111000001101101110010",
    804 => "01111110111111111010111001001001",
    805 => "01110101111111111011100101010011",
    806 => "11011111111111111110000100011001",
    807 => "01101111111110110110111100001111",
    808 => "11110111111011110011101001101000",
    809 => "01011111101111110111001011000010",
    810 => "10111111100000000000000000000000",
    811 => "11111010101011111110010011011001",
    812 => "01000111011101110010100000000000",
    813 => "01111010100110011011101100111111",
    814 => "01011101110001101101001100100001",
    815 => "11111111011111100100010001110010",
    816 => "11001100111110111000111001000001",
    817 => "01100100011101110000010001100001",
    818 => "11111101101101100001000000100001",
    819 => "11110001001111110101001000000000",
    820 => "11110001011011110101010100110010",
    821 => "11011111111111100101010100011101",
    822 => "11101111110111111001100011110001",
    823 => "10111111100000000000000000000000",
    824 => "01111111011111000101010100101101",
    825 => "01111100110101111110110010001111",
    826 => "11101111110011111000000001100111",
    827 => "01011011101111011100011101011010",
    828 => "00111111100000000000000000000000",
    829 => "10111111100000000000000000000000",
    830 => "11011011101100111101100010101101",
    831 => "11011101000111100011110110001000",
    832 => "01001111111010010001001010110011",
    833 => "01100110101110111001101011000010",
    834 => "11101111111101110011111011100100",
    835 => "10111111100000000000000000000000",
    836 => "11111011101011110111001110001010",
    837 => "01111001111110011110101100010101",
    838 => "01111011011111010000010011111011",
    839 => "11011110110111011111100110000110",
    840 => "11111111010111111011111100000110",
    841 => "10111111100000000000000000000000",
    842 => "11010101111101111101001010110000",
    843 => "11111111011110111000110111011101",
    844 => "01101000111000000001111000100001",
    845 => "01111101101001110100101000010110",
    846 => "11011011001101101111000100000111",
    847 => "01011100111011010010111010001011",
    848 => "10111111100000000000000000000000",
    849 => "11101011000011010100101001001111",
    850 => "01001111111010110111000111001111",
    851 => "11111011111001110110101001110000",
    852 => "11101110010101011010010010010000",
    853 => "01111011111000100100100011111110",
    854 => "10111111100000000000000000000000",
    855 => "10111111100000000000000000000000",
    856 => "11100011111100111110011011001011",
    857 => "01111000101110110110110111110100",
    858 => "11010110111111101110111111001101",
    859 => "01111110011101011101011000001111",
    860 => "11111101110111101111111100101110",
    861 => "10111111100000000000000000000000",
    862 => "11111001100111111100111111011110",
    863 => "11011111111000101101011000101011",
    864 => "01111011001110111110010110010001",
    865 => "01101111111011111011000100111100",
    866 => "01110110110111101010010011011011",
    867 => "11111100101000100110100010010101",
    868 => "01010101001000110111011101010111",
    869 => "01011111111101110111010001101010",
    870 => "11111010010111111110000110100011",
    871 => "11111011111100001011011010111101",
    872 => "01111011101011111010010011011100",
    873 => "11011101100110111010100100010000",
    874 => "01011101111111111100111001101010",
    875 => "11111011111111011100111111101010",
    876 => "11011111011101111000011100101110",
    877 => "01111101101010111110001010001011",
    878 => "01001011001011001011011111110101",
    879 => "11110110111111011101110010101100",
    880 => "01010101110101110011101010100100",
    881 => "11111111001111101110010000000001",
    882 => "11100101111101001011001000100101",
    883 => "01101101111011111001000101101100",
    884 => "11011100111011011011000100110100",
    885 => "11001111110011110110000101110011",
    886 => "01101111110111010100101000100110",
    887 => "00111111100000000000000000000000",
    888 => "10111111100000000000000000000000",
    889 => "01111011101011011101100011110100",
    890 => "11000000000000000000000000000000",
    891 => "01101101101010111111011000001110",
    892 => "11111011100111110000100110100011",
    893 => "11111110111101111001111110110100",
    894 => "00111111100000000000000000000000",
    895 => "01111100111110001010101010111011",
    896 => "11111010101111111001010011011110",
    897 => "11110111111101011000100111011110",
    898 => "11010111010111001100101010000001",
    899 => "11111110011111010010011000101111",
    900 => "01001010101111001110111000010100",
    901 => "11001101011111011001110100101000",
    902 => "01111111011111111101000001101101",
    903 => "11111101111100111101110001111001",
    904 => "11011011101111110010101110111100",
    905 => "01101101111101111010110010010111",
    906 => "01001110011011111111000100100111",
    907 => "01111000111110111000001100010100",
    908 => "01111101110011110001111000010000",
    909 => "11000000000000000000000000000000",
    910 => "01111110111111110010100010001001",
    911 => "11111011000110111010100101000000",
    912 => "11101111111111110100101011100110",
    913 => "10111111100000000000000000000000",
    914 => "11101111111011111100001001001000",
    915 => "10111111100000000000000000000000",
    916 => "01111101111000000101011110100110",
    917 => "01001001110111111110001101001000",
    918 => "10111111100000000000000000000000",
    919 => "11111111001111110101111010100001",
    920 => "01111110111110010001001000100011",
    921 => "01110011100110110010111110011111",
    922 => "11111011111111110111011000001000",
    923 => "11101100111111100011011010100010",
    924 => "10111111100000000000000000000000",
    925 => "10111111100000000000000000000000",
    926 => "11011000111101110010101110101011",
    927 => "10111111100000000000000000000000",
    928 => "11011101111111111011001100101100",
    929 => "01010111110011001110101000011110",
    930 => "01110100010010100101001110100000",
    931 => "10111111100000000000000000000000",
    932 => "01011101100111000010111011110010",
    933 => "01111110101110101111111101001010",
    934 => "01110101010101111010000000110000",
    935 => "11011110111111100011011101110001",
    936 => "11011111111011010011011001000001",
    937 => "11001011111101110110000110000110",
    938 => "10111111100000000000000000000000",
    939 => "01011111110100110001101111111001",
    940 => "11011111111011110100010010110100",
    941 => "11110110111111110001001110010000",
    942 => "11111101101111111101100111111000",
    943 => "11111000111010110101000111111001",
    944 => "10111111100000000000000000000000",
    945 => "01011110111111111111100100001111",
    946 => "11111010011110111111000000011011",
    947 => "11111001010110110110110101011110",
    948 => "10111111100000000000000000000000",
    949 => "11101011111111110110011100011110",
    950 => "11100110001111101101010000011001",
    951 => "11110110011111111110001011101111",
    952 => "01111111011110111100111000001110",
    953 => "11111110111001100110111000100110",
    954 => "01111011001101100001100100001001",
    955 => "01101111110101111101010110011110",
    956 => "10111111100000000000000000000000",
    957 => "01111011011011101111111010000101",
    958 => "01111011101000110110001101100110",
    959 => "11011011000111110111111011101011",
    960 => "11111110001011011101011001110011",
    961 => "01001011000110110011110111100011",
    962 => "10111111100000000000000000000000",
    963 => "01010001011111110001111110111011",
    964 => "11101111110011010110110001011011",
    965 => "11111010100110100010110010110110",
    966 => "01110111101111111001010111001111",
    967 => "01111111011111110101001110010100",
    968 => "11100101101100111011000011000010",
    969 => "11111111011001110010000011100110",
    970 => "11110101101011110011000010011110",
    971 => "10111111100000000000000000000000",
    972 => "00111111100000000000000000000000",
    973 => "11011110011111110000001011011100",
    974 => "01100100111111110100100001000101",
    975 => "10111111100000000000000000000000",
    976 => "10111111100000000000000000000000",
    977 => "11101011100110110011111000011110",
    978 => "01101010111101010110111100010110",
    979 => "11011011111110011011000010010011",
    980 => "01110101111101110111000001010010",
    981 => "10111111100000000000000000000000",
    982 => "11101110111111100001000010011100",
    983 => "11000000000000000000000000000000",
    984 => "10111111100000000000000000000000",
    985 => "11100111011111111100101101010110",
    986 => "11101110001110110111101001110100",
    987 => "11000111101111011010001000000000",
    988 => "11011100110010110000111011110001",
    989 => "01110101100001110100110000011000",
    990 => "10111111100000000000000000000000",
    991 => "01101111111011111111000111010000",
    992 => "01111000111111110011001111110011",
    993 => "11111011111110001001101001110111",
    994 => "01011111011011110110010111001011",
    995 => "11111110101111101001000011000001",
    996 => "01101110110111111010110001100000",
    997 => "11111101111111010110011101010110",
    998 => "11011101111110101111110011100100",
    999 => "11111111011001000010011011000011");


  component floor is
    port (A : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          Q : out std_logic_vector (31 downto 0));
  end component floor;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (3 downto 0) of std_logic_vector (31 downto 0);
  signal cc : std_logic_vector (31 downto 0) := (others => '0');  
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
begin  -- architecture floor_tb

  i_floor : floor port map (s_a,clk,c);

  judge: process (clk) is
  begin  -- process judge
    if rising_edge (clk) then  -- rising clock edge
      ccc <= cc ;
      if ccc = c then
        Q <= x"30";
      else
        Q <= x"31";
      end if;
    end if;
  end process judge;

  ram_loop: process (clk) is
    variable ss : character;

  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      s_a <= a_lut (addr);
      cc <= ans_lut (addr);      
      if addr >= 999 then
        addr <= 0;
      else
        addr <= addr + 1;
      end if;
    end if;
  end process ram_loop;

end architecture;
