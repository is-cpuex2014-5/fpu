library  ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity fneg_tb is  
  port (
    clk : in std_logic;
    isRunning : out std_logic;
    result : out std_logic);
end entity fneg_tb;

architecture testbench of fneg_tb is
  constant array_max : integer := 999;
  type lut is array ( 0 to array_max) of std_logic_vector(31 downto 0);
  constant a_lut : lut := (
    0 => "01101111111101010111011101101110",
    1 => "01011111011111011011001010010100",
    2 => "01011101101111111001011101101001",
    3 => "11111101111101111101011111110011",
    4 => "11101110101111111011100101011101",
    5 => "00101010101111110011010111011000",
    6 => "00010011101110110001110111110101",
    7 => "01001100111101100011010011001000",
    8 => "11111101010111111010011100000000",
    9 => "11111011011111110100111010110111",
    10 => "11111011110111010010111000111000",
    11 => "11101111100111111111111111011011",
    12 => "00110111100111110100111001001010",
    13 => "11011011011111010111010001111111",
    14 => "11110111111111110001101111001010",
    15 => "11011111101110110101000010100010",
    16 => "00010111001111100011011010000110",
    17 => "11101101111111111110110101010101",
    18 => "11000111010111100101100011010011",
    19 => "01010110101110101000011101110000",
    20 => "11011101011110110011110001100001",
    21 => "01110111001010011101000011101010",
    22 => "01110111111111110000111001001100",
    23 => "01111101100101110000010110000011",
    24 => "01110111111110110101000010011100",
    25 => "10011111111011111101100011010001",
    26 => "01101101110110011000011000000101",
    27 => "10110101110101100111101001100011",
    28 => "11001011111101010001010000110101",
    29 => "01101011101111110011010100001001",
    30 => "00111011011111101100111000111100",
    31 => "00100111011111110001100010101010",
    32 => "11111000101110111110011110100110",
    33 => "11111111010110110011100101000000",
    34 => "01110101111011010101110101100010",
    35 => "01101110011011100101010001100100",
    36 => "01101011101100111110011011001010",
    37 => "00101101010110111011111110110011",
    38 => "01011111110011110010000000001001",
    39 => "11111100110111100110110000111011",
    40 => "11111110111011111010111100110110",
    41 => "01101111111111110100011000101010",
    42 => "11101111001111111111010010011111",
    43 => "11011110110110111010010100011010",
    44 => "11111101110111101110101101111000",
    45 => "11110011010111111110100111101010",
    46 => "00101011101010110101110111011110",
    47 => "10110111101011111001100011001011",
    48 => "10001111110000110001100100111101",
    49 => "11111000111110110110101111100011",
    50 => "11101011111111001001100100001110",
    51 => "01010111110110111110100101000000",
    52 => "10011111011101101000010011000110",
    53 => "11011110111110111111011110001011",
    54 => "11001011111111111100001000010000",
    55 => "11111110101111110010010101010000",
    56 => "11011011011010110101010010110110",
    57 => "01000110111111100111100110001010",
    58 => "01101111111111011000100000101111",
    59 => "11100111011011110001001101001100",
    60 => "01111101111101011000011010011111",
    61 => "00011111111011101010000101001110",
    62 => "10111011111110110010110000000001",
    63 => "01110111111111111001111100000000",
    64 => "01011010111001000001101010011110",
    65 => "11110011101111000001111000110000",
    66 => "01100111011100111001011011010000",
    67 => "01011111100111111011100011110110",
    68 => "11110010111010111001111111100111",
    69 => "01101011111111111110011010001000",
    70 => "00111111110110100011110000011101",
    71 => "11111011110110110001100010100110",
    72 => "10110110101111111101011001000011",
    73 => "01011111011101111101000100000001",
    74 => "11111101010111111111010110100100",
    75 => "01111101010111110100010010000001",
    76 => "11101101110011110101100111000010",
    77 => "10111111111010111001101110101110",
    78 => "00111110111111110111000010101010",
    79 => "10001011111110001100101100000010",
    80 => "11111011001101100100010110010010",
    81 => "11011110011100110011111011110101",
    82 => "11111100110011111111011111111010",
    83 => "11011111100111101010100001101101",
    84 => "11100100110010111111001010000001",
    85 => "01001011001111111110101001011010",
    86 => "11000110110111100111010101011110",
    87 => "01100111011111111001110101010111",
    88 => "10111010111111110001111100010001",
    89 => "01101111110111110010101010101101",
    90 => "11010110011111110000111100111111",
    91 => "10101010111111010100100101100001",
    92 => "11111011100111000000101000110010",
    93 => "01111011111011110100010101010100",
    94 => "11100100010110011011111001100111",
    95 => "10101111001111100000011110010001",
    96 => "00100101111110110011111110010100",
    97 => "01111010011101011101111000001101",
    98 => "11101110111101110000100100101100",
    99 => "11011111111100111000100100000101",
    100 => "10111101101111111100010011101010",
    101 => "01111101110111110000101110101000",
    102 => "01110111000011110111010000000110",
    103 => "01111110011111100010011110111011",
    104 => "00101111011111110000111100010110",
    105 => "01111110111010100101001101101101",
    106 => "01011001110101010011100010000100",
    107 => "01100101001101111101100010110100",
    108 => "01110100111111111100000011011111",
    109 => "01100010011111000011111110100000",
    110 => "01011101111111110111100110001011",
    111 => "11111110111101110011001010001001",
    112 => "11001111101111100100101001011001",
    113 => "01111110111111011011010111000011",
    114 => "01011101011101110111011111100011",
    115 => "10100110111110111010100000000001",
    116 => "11111011011111110110100111001000",
    117 => "10100011110011111101101101100100",
    118 => "11111100000111100000110101000100",
    119 => "11011111011011111110001001100010",
    120 => "00100011101011110000100100000001",
    121 => "11110011101011101100111010010111",
    122 => "00000011011110110011111110110000",
    123 => "00110101111001010000010101000011",
    124 => "00000110100001110111000011100111",
    125 => "10111011110100111001010011011111",
    126 => "10111111110100001100110010110001",
    127 => "10000111111101110111001100101001",
    128 => "11101111111111111100111011101010",
    129 => "01011111111111011010110000111101",
    130 => "01010111001111110000010001010001",
    131 => "01111110011110011100110111000111",
    132 => "10111011111110110100111110101110",
    133 => "01111110111111110001000001100101",
    134 => "11110011111001110101110101000011",
    135 => "01111111011111000010101100010101",
    136 => "01010110111110111110100011010000",
    137 => "11101110101100111111101011001110",
    138 => "01101011101101010111101000111111",
    139 => "00111111100111111111010010011001",
    140 => "11010001010111100010011011110101",
    141 => "10111011001111101011101100101111",
    142 => "10111110100110110100001110111111",
    143 => "11101111111111100100000111111110",
    144 => "01100111011011111101000011100110",
    145 => "10011110101011010100010000111011",
    146 => "10111011111110011011010001101000",
    147 => "11010100110111110100011111011000",
    148 => "10110111110110111111000011011011",
    149 => "01011011111101011011011110010101",
    150 => "11011100010111110000101101011111",
    151 => "11111110001011110001010110011110",
    152 => "00111010011011110010000011011001",
    153 => "10011011101110101110001001000011",
    154 => "11110111111111100111110000100001",
    155 => "10100011011101111010101000110110",
    156 => "01100111111011111001100000100110",
    157 => "11011111111011110011110100110101",
    158 => "01111111001101111110111101111110",
    159 => "11001111011011011100101111100010",
    160 => "00110011100111111100010110000010",
    161 => "10111110111011111010010000000111",
    162 => "11111100111001110011111010110111",
    163 => "11110111110111110100110000000110",
    164 => "11101111111101111100001010101011",
    165 => "11101111111101010100101110010101",
    166 => "00101101111110001101011011011101",
    167 => "01111110111111110111111010011100",
    168 => "00111000110110110000010010110100",
    169 => "10111101110110111111011000010101",
    170 => "01010110111110101011001001111101",
    171 => "01110111111111110011111000011100",
    172 => "10111111111111110101010011000000",
    173 => "11111010111111111111000111101001",
    174 => "00110111111111110100010000011001",
    175 => "10110111111111101000110110101001",
    176 => "00111110011111110010011011101101",
    177 => "11101111101110111110011110000110",
    178 => "01111111010110110000010011101110",
    179 => "11011011110011001100110100011101",
    180 => "01001111111110010110000011110100",
    181 => "01101101101011110010111011001010",
    182 => "01101110111111110111010010001100",
    183 => "00001010101001101000000001111100",
    184 => "11111110111111011011111111100110",
    185 => "01011111111101111000001010100101",
    186 => "01110101110011110101101111000110",
    187 => "11011111111101100000110101101101",
    188 => "10011011100111111010010100101111",
    189 => "11101100101111010011000000000000",
    190 => "01010111111011101101100110010100",
    191 => "11111110110110101011010110110100",
    192 => "10011011111110110100101010100001",
    193 => "10101011111101111011101001001110",
    194 => "11111101011110111100111010001011",
    195 => "01011111011111110001000100111110",
    196 => "00111011110100110000110111111000",
    197 => "01111111011101100100010111011100",
    198 => "11010111110110101000111100000101",
    199 => "01101110111011110111000011001000",
    200 => "11111011111011111000010011110000",
    201 => "11100101111101110110001110010010",
    202 => "01111111001010111000000010010111",
    203 => "10110111110101110000110000010111",
    204 => "11110111111110111101100101000111",
    205 => "11101110111111111100100000011101",
    206 => "00111011111111101100010000101101",
    207 => "11111111011111011011111001010100",
    208 => "11011111101101110110011110010101",
    209 => "01110101100111110010001101110000",
    210 => "01111111010111001110001101010011",
    211 => "01110011111111111101101110101111",
    212 => "01011110111110000010111110100101",
    213 => "11111110100101111100000101000101",
    214 => "01101110110111110011111111100110",
    215 => "10101111111111101001010101001100",
    216 => "01011111111110111001010111010111",
    217 => "10101011111111101011010100001110",
    218 => "10111110110101111100011001111010",
    219 => "01001111111101110001110101010001",
    220 => "00111111001111111010000101010110",
    221 => "00111111110111010000111101110111",
    222 => "00110111111001110010111100111100",
    223 => "01010011100011111010011101100101",
    224 => "11011011011101011001110000110100",
    225 => "01110111011111011100111110001101",
    226 => "01001111011101111000000001101110",
    227 => "00111111111110110110101100000101",
    228 => "01110111110111111011011101010101",
    229 => "11111011011111111010001011001011",
    230 => "01101010111111001111101010111001",
    231 => "00011111101010111000000010110000",
    232 => "00111011101001100111011000101011",
    233 => "01010011111111110100011100101001",
    234 => "01110111101100011000000110110000",
    235 => "11111110111011110111001001000110",
    236 => "00011001111011101000100110001000",
    237 => "00110111111111011100001101111100",
    238 => "01111110111001011001110011000001",
    239 => "01111101111111111111000110010101",
    240 => "01110110000111101000111010010010",
    241 => "11111001111101110111101111000001",
    242 => "00110111100111111000011110111111",
    243 => "10111111010111011111101001110011",
    244 => "11011111011111101001111101111010",
    245 => "10011010101101111010010101110110",
    246 => "00110111011101111100011110100011",
    247 => "11111001011101110100100000101101",
    248 => "11011001111111100111111000111101",
    249 => "11111110101101110101000000001000",
    250 => "11111001111101110111101011001010",
    251 => "00111111010111110000101000101111",
    252 => "10111110111101011111111101001101",
    253 => "11111001111111111000011010101011",
    254 => "00011111001111110001001100111110",
    255 => "10001110111111110110001011100110",
    256 => "11101111101001010000111011010100",
    257 => "01101011111001111100001000010110",
    258 => "01101101110110101001111000000011",
    259 => "01011111111110111010011010000110",
    260 => "01101110011110011111101111000011",
    261 => "11101110110010010110100110100000",
    262 => "11111101110111101010101111110111",
    263 => "00101110011101101010011101100111",
    264 => "11110111011011110111101110101100",
    265 => "11111110111111110001101010111000",
    266 => "00110101111111111101000100000000",
    267 => "11010101010111110011010010111101",
    268 => "11011111001111111100000100101111",
    269 => "01101110101101101101000010100101",
    270 => "00111011111111000000111010111011",
    271 => "11111100101111101110100011000000",
    272 => "10101111110101111001000110111100",
    273 => "11111101011111111111000000111000",
    274 => "11101110111111110000101110100110",
    275 => "11111111010111101101001110011011",
    276 => "11101011110111110111110111001001",
    277 => "11111110100111100001001100111011",
    278 => "11011111001110110111101110100011",
    279 => "00111110111110111011111000101001",
    280 => "00111110111111110101110001101011",
    281 => "11101111001001110001110001100011",
    282 => "01101101111111111001011000010011",
    283 => "10111011101110100111101110100110",
    284 => "10110111011011100110011001110011",
    285 => "01110111000111100011110011101001",
    286 => "00010100100101011001101000001101",
    287 => "01110100011000111111100101101100",
    288 => "01110111111111111111111011011000",
    289 => "01110011001110110001111110111010",
    290 => "11011111111111010010100110111011",
    291 => "10010111111110111111000100100110",
    292 => "11101111111110011101100000110000",
    293 => "01111011010110011101011000111100",
    294 => "11111100110110101101101110001111",
    295 => "00111111111110111010100010111110",
    296 => "11101101001111011111101100010101",
    297 => "11111101111111110010011000100010",
    298 => "10111011111111011101000110111100",
    299 => "01111010011011110010010010101010",
    300 => "01111001100111010101100011101111",
    301 => "11111011111111101010101001001001",
    302 => "10100111111111110111001000011001",
    303 => "10001111100111110001101011101011",
    304 => "01111110111011111000001100000101",
    305 => "01111110011010110010001001110111",
    306 => "11111110111001111101110001010000",
    307 => "11111011110011010010001101111011",
    308 => "11111111011110110011001111000001",
    309 => "10101111111011110011011100000110",
    310 => "01011101001110001010000110100000",
    311 => "01111011110111000011001100010010",
    312 => "01010111101111111111111011110001",
    313 => "01010111111101001010101110001011",
    314 => "01010111110111011011100101010001",
    315 => "01101011011010100100101011011100",
    316 => "11111010011111001111100110001011",
    317 => "00110110011111101001110001011011",
    318 => "00111111011001100011100101010101",
    319 => "01111011111111100101100100011101",
    320 => "00111101011011111001001110001100",
    321 => "10011011011101111110011111111011",
    322 => "10111110111100001011011000010010",
    323 => "11101111100111110110011010110100",
    324 => "00101001011111100011000010111011",
    325 => "01100111111011110100101001000001",
    326 => "01001111001111110111101110110000",
    327 => "01110111001111111011101110001010",
    328 => "01110111111110111010000100010011",
    329 => "11111011111011110111110100010000",
    330 => "01110110101111111010000001000101",
    331 => "00111100101101111001111000101011",
    332 => "11011111101010011000101100010010",
    333 => "11101111101111110101110000000001",
    334 => "11101111101011110011001101001101",
    335 => "01011101111111111010011010010101",
    336 => "01111110111001110001001111110110",
    337 => "01111011111110101001000001101001",
    338 => "11000101011111100100100111000000",
    339 => "11011101100101011000001011111110",
    340 => "11111110101011110010010011110001",
    341 => "11110110111111101101110100110011",
    342 => "01111110111001110010010111101010",
    343 => "11110111111110110101010101010111",
    344 => "11110101101111110110101000110110",
    345 => "01001010111101010001100110010110",
    346 => "11110110101110110011001000111110",
    347 => "10011110011111111101111111100010",
    348 => "01011011011101101000100011010111",
    349 => "11101110011101010111110111001101",
    350 => "11110011111010011010010000001101",
    351 => "01110100111101111000000100001001",
    352 => "11011011111011010010101110010010",
    353 => "10111110111100011111010110011010",
    354 => "01011110111011000101111011001010",
    355 => "11011111001110111111101100001000",
    356 => "01011010110111111011101001000100",
    357 => "01101100111110100111011000100100",
    358 => "11101111101111100100010111111100",
    359 => "01111000001111110010110011011100",
    360 => "00011110111111100011010001100010",
    361 => "11111110011101110001111111101110",
    362 => "11111100111110110101111110101110",
    363 => "01100111111111111010100010101001",
    364 => "01101011101110110110110111001000",
    365 => "11111011011110110011100000110010",
    366 => "01110011110011110100011111101011",
    367 => "11110111001111110100100001011001",
    368 => "01110011111000011000111101000100",
    369 => "01001001111111111100100001010100",
    370 => "00111110011111111001001111000000",
    371 => "11111001101111110110111000000011",
    372 => "10111111111111111100111000110010",
    373 => "01100111100111110101000111110111",
    374 => "01011110011111111010011110011110",
    375 => "00011111011111101101110010111000",
    376 => "11010111011001111000010001101100",
    377 => "11110010111101010010001100111000",
    378 => "01011111111110111010111100010100",
    379 => "11100011110110101000101110001111",
    380 => "11010011011110101000100100111000",
    381 => "11010111100101011111011011010110",
    382 => "11110111011110111100100010100101",
    383 => "10110000111110110001010011110010",
    384 => "10101001101110101100111110100100",
    385 => "10111101111101111000001001101111",
    386 => "11010101011101111101100010000111",
    387 => "11101100001001011010000000111001",
    388 => "01101111001111110010110011011000",
    389 => "00001001101101010100011110110001",
    390 => "11111100000111100111111110000100",
    391 => "11101111111111111000111011110010",
    392 => "00111110100011101011111001010010",
    393 => "10011111111111111110000110010110",
    394 => "11011011111011010001110101011100",
    395 => "11100110010000010101100011110000",
    396 => "00101111111011000111011011111011",
    397 => "01110111111011110001011010010101",
    398 => "10011011100101000110101111010011",
    399 => "01011111010110111110010000010011",
    400 => "10000110010011110110110101101011",
    401 => "11111110011001001100010001111111",
    402 => "00111100111110011110010001010100",
    403 => "01110011110111101010001111010101",
    404 => "01111010110101111101100001001111",
    405 => "11010111111111010000011010010100",
    406 => "01101101101111010111000011001110",
    407 => "01111111011111001110000010000011",
    408 => "11111101000111110010101011010001",
    409 => "11001011111110011110001111100000",
    410 => "01101011100010111011011110000101",
    411 => "01101011111110111010000101001010",
    412 => "10001101110111010000001010001000",
    413 => "01111101001100110000100110101001",
    414 => "11101111111111110000101000110111",
    415 => "11101111101011100011100001100100",
    416 => "00011111101110110101000111010101",
    417 => "01011010111111101110000011010100",
    418 => "01110101111000101010011101010100",
    419 => "10011111111101110101110100100110",
    420 => "11111001110100011010010000000110",
    421 => "11111110110110011000010110110110",
    422 => "01111001101101111100111001001101",
    423 => "00100111011111000101100000110001",
    424 => "00011111111101111100010001110011",
    425 => "01100101111111111000101010111111",
    426 => "10011101010001110011001100010000",
    427 => "11011110110101111110101100011010",
    428 => "11110100110001111111110100111011",
    429 => "01001111111100111100011011110110",
    430 => "11111111010110101110001011000001",
    431 => "01110101100111111011010101111111",
    432 => "10110111110111110001000000001101",
    433 => "11110111011000111000110100000000",
    434 => "11101110001011101110011111110101",
    435 => "11001111111111110011111100111001",
    436 => "11010111111101101101001101101000",
    437 => "10100001111111010101101011010011",
    438 => "10110011110111110010111010000111",
    439 => "11110110111110101100001011110001",
    440 => "01011111101110111100001010111100",
    441 => "11111101110011100101100010110111",
    442 => "01110111110100111101101011111000",
    443 => "11111100011100111001000010001111",
    444 => "01011111111111110011100010010100",
    445 => "10010111011101010101011011100000",
    446 => "01100110111011100100111111101100",
    447 => "11011110111111010010101101111000",
    448 => "01010111111111110001111001010000",
    449 => "01011111111010111100011100010011",
    450 => "11111011011111111001111101101000",
    451 => "11111110011111100010001001111001",
    452 => "01010011000110000011110000110000",
    453 => "11111111001110111010110101000001",
    454 => "11111100101110010100110011010011",
    455 => "00111111111111110110010111001001",
    456 => "11110111010111011110000010000010",
    457 => "00011001110101111111111111111111",
    458 => "11011111111001110100110111011110",
    459 => "10100100111111110011010001101100",
    460 => "11010100111110010111010011001010",
    461 => "11111101010110100000101110101101",
    462 => "01101110010110101011001110101111",
    463 => "01010111110111111000011110000110",
    464 => "10111011000001011100001011010011",
    465 => "00111111111110111111111000100101",
    466 => "01101011111111110110101010010001",
    467 => "11111011010110111101101110101100",
    468 => "10111110111111110111001011000100",
    469 => "01110010110100111100011010110011",
    470 => "00011100100110011101010101000110",
    471 => "01001011111101110101001001101000",
    472 => "11100111111110111011100101010000",
    473 => "11010101111111011000111000001011",
    474 => "11101111111111010110011101110100",
    475 => "01111111011100111110111011111010",
    476 => "01110111101001110001011110101000",
    477 => "11011111011111110110111000111010",
    478 => "00111111110010111101100101111110",
    479 => "11010111111011011011011000100010",
    480 => "01110110111101010101101001111100",
    481 => "00111111101011110010001010011100",
    482 => "11010111111000111111000100001110",
    483 => "10110111110000111111001001011000",
    484 => "11011111111111110000100000100011",
    485 => "01011110110010111100110001010011",
    486 => "11101101111111111101000101010000",
    487 => "01111111011110110010000110111101",
    488 => "11011111011110110100101010100001",
    489 => "00111111100110110100111010101011",
    490 => "01110110111110111010010001010100",
    491 => "00010010101011111011000000011100",
    492 => "11111100111111110100000011001110",
    493 => "00111111010111011100111000011101",
    494 => "10000100111111111110110000011111",
    495 => "01000111110111111111000111110001",
    496 => "00011111101011111010010011110011",
    497 => "10011111100101100111110011000100",
    498 => "01101111001111111010100111101110",
    499 => "10110011100110010100110111000011",
    500 => "00011011101101110011011010111010",
    501 => "00001010011110110000110010011101",
    502 => "01111110010110101001111110111010",
    503 => "11111010010110110110011101100110",
    504 => "10110110011111101011011110001100",
    505 => "01011011111100010010001111110110",
    506 => "11011101110111110001110001100101",
    507 => "01111101001101110110111001101111",
    508 => "00111110110111011010010010110000",
    509 => "11110000110011110111011110000001",
    510 => "01101111111111111101011101101011",
    511 => "01010101111011110111110111111111",
    512 => "01011111100001111100001101001100",
    513 => "11110111100111100110001110011011",
    514 => "01010111111111110000001000010001",
    515 => "01111001111111010001010011110110",
    516 => "11001110101010101110110110110000",
    517 => "01010101101011110001111110001010",
    518 => "10110111111110111110010110111010",
    519 => "10111110011110101001100100100011",
    520 => "01110110111111101101001101011111",
    521 => "11010101001111110001101100111010",
    522 => "11111011101001010111101000010110",
    523 => "11111001010111111111100111101010",
    524 => "11110101111111010100011011010100",
    525 => "01011011001100110010000000000011",
    526 => "11111010010110110011111100110001",
    527 => "11111010111111000000010000100111",
    528 => "01000110111111011110000010011110",
    529 => "11111101100111111010011000100010",
    530 => "11011111110111100110111110110000",
    531 => "11011111111111101100001000010111",
    532 => "11111110011111111010010101111001",
    533 => "11101011001101111100101100101010",
    534 => "01101101010011011000000101001101",
    535 => "01010110101011110001010110011110",
    536 => "00111001110111010111010011110010",
    537 => "11111111011010001110100011010111",
    538 => "11100011111011010010001101111101",
    539 => "01101111011100111110011100011110",
    540 => "00110111111000101101100001101101",
    541 => "00010111111111110111010001110010",
    542 => "01111011100111110000000100100100",
    543 => "11111011110100111011101001101011",
    544 => "01101100110011010111111011010001",
    545 => "11111110100101101101011101011000",
    546 => "10011111011111111111010001011111",
    547 => "11011101110110110111110110111100",
    548 => "01001101111011111000001111101010",
    549 => "00000111001101110010010100001100",
    550 => "01111011111110111010110100110100",
    551 => "00111110111001110101100111100011",
    552 => "01000110101111100110101110000010",
    553 => "11011110111111110001000100101110",
    554 => "11111101010011010010010101111011",
    555 => "01111101111011111111111101101111",
    556 => "00101010111101110001010110000111",
    557 => "11001111111101101110011001011100",
    558 => "01100111001011011110001001010110",
    559 => "11111101101011100011000001111111",
    560 => "00100110110111110101001110101111",
    561 => "11110001011111100101001100011110",
    562 => "11110111000011111011111010111000",
    563 => "11100011110111000001101001010010",
    564 => "11010111101011111101110000111111",
    565 => "01111110001101110001111001101111",
    566 => "11101101111110011110100110101100",
    567 => "11111010111110110111100011011100",
    568 => "11111110111111110001100011110001",
    569 => "01011111011101101111001100101000",
    570 => "11110111101111111001110001000000",
    571 => "10111001110110111000000000000101",
    572 => "01101110111111011111001100101010",
    573 => "11110111100010111000000110111010",
    574 => "10110011011110111100101110001110",
    575 => "00011111101111111000111100101111",
    576 => "11110111010111111101011100011001",
    577 => "11111101111110011111000010101010",
    578 => "01101010111111111011100101010101",
    579 => "11011111111111110111100110010101",
    580 => "10011000111001111101001010000011",
    581 => "11111111011111111100101110110110",
    582 => "01100111111100100010000111110110",
    583 => "00111011111011111011011100001010",
    584 => "11101111001101101110001011101010",
    585 => "11011101011011101001110011001001",
    586 => "11101111111111000011000011110010",
    587 => "10110011111111010011001110001111",
    588 => "11111111010111010110010101110101",
    589 => "11110110101001110110010011100111",
    590 => "00111110110011100001111001011011",
    591 => "00001111111101011101011011110010",
    592 => "10110110111001111101000111010001",
    593 => "01101011011111100001101000000010",
    594 => "11111100111001110010010111011100",
    595 => "11110101111100101110001101101011",
    596 => "00011101111110111010100010110100",
    597 => "01011111101111110011011000100101",
    598 => "01011011011011110100000001001000",
    599 => "11011111111101110000100111110001",
    600 => "10101110111111111001100000111001",
    601 => "11011101101111110101101010011111",
    602 => "10001111011111110011011010101111",
    603 => "10011111011111010111101111011001",
    604 => "11100011110001011000110101001011",
    605 => "10101011101101111001000011001000",
    606 => "11101111100110111011101010101100",
    607 => "11111101101111101111100000000010",
    608 => "01011111111111100011100111110111",
    609 => "00011111011100111100000100110011",
    610 => "01101001111010100000111101110000",
    611 => "01000111111111010010001011000011",
    612 => "01110011111110111100100110100111",
    613 => "11111011100111010101111010100100",
    614 => "11111110110111101111000001111100",
    615 => "10110111011100101100000000001010",
    616 => "00111111111001111101100101001001",
    617 => "01101111100111010100110100100110",
    618 => "01111101011111110001001000111100",
    619 => "11101100111111100100010110101001",
    620 => "00111101101110110010011111110100",
    621 => "01100111111110111010000110010111",
    622 => "01111010110110110101101110001001",
    623 => "01101010111110110111111101001110",
    624 => "10101110100100111100110010110010",
    625 => "10010111110110011011000010001111",
    626 => "00001111001101010000010100011101",
    627 => "11100100111101110000011000010010",
    628 => "11111110110111100100000010110101",
    629 => "01111011111111111001010101001000",
    630 => "11110010111111100000000111111111",
    631 => "01111110101000111000000010010011",
    632 => "10110011111111111100000001011101",
    633 => "00011110100011110101100000000101",
    634 => "01011011010111110100001110110010",
    635 => "10011111001111111110000111100100",
    636 => "01101001101100100110010000011001",
    637 => "01110100111011100000101000110110",
    638 => "11111011111001110000001101000100",
    639 => "01111100111010111100011100100101",
    640 => "01111001111101111100100111111001",
    641 => "11010101111111111111110111111010",
    642 => "01111110101111110001010101011101",
    643 => "10111011101111111001011000100111",
    644 => "10011010011001100101100010101110",
    645 => "11011111010010011000110100010011",
    646 => "01101111110011010110110000010001",
    647 => "11001011111011110101001101111000",
    648 => "10111111011011111000111011000110",
    649 => "01111001101110111100110100011000",
    650 => "01111111001101010011011001100110",
    651 => "01101001110111001101000111011101",
    652 => "11010111111010110110000111111101",
    653 => "00111101001110111111101101100010",
    654 => "11100111010111111101110110000010",
    655 => "00101111111011100001101000101100",
    656 => "01111010110110100001101000111100",
    657 => "10111111010111001100001110110101",
    658 => "11111010011011011111010011000001",
    659 => "01111010011111011000100101001011",
    660 => "00011010110110011000001111110110",
    661 => "01110111101111101101111101100011",
    662 => "01011101110011101000100010111100",
    663 => "01011111110110101000001000111111",
    664 => "11101100111111010101011001100110",
    665 => "01110101110011010010111110111011",
    666 => "00001101011111110000110101100000",
    667 => "01101111111110100001011100100100",
    668 => "11111100100011111110100010111011",
    669 => "00101111111101111101011100110010",
    670 => "11110001111111101101100000011001",
    671 => "10011111111011110111010111000010",
    672 => "11011001110111101001100010111110",
    673 => "11011101111111110001011001001100",
    674 => "10111111100111110111101000001011",
    675 => "11111110011111011101010110111000",
    676 => "10111111001111011011011110101000",
    677 => "01000110011011010100111100001111",
    678 => "11011101010111101100101011100110",
    679 => "01100101111111111001101011111111",
    680 => "11011010111111111011010110001011",
    681 => "11011010111010110111001100010101",
    682 => "10011111101110011101011111111000",
    683 => "11001000101111110010101010000110",
    684 => "01001011101110100011011011000100",
    685 => "01011110111111011100001110011011",
    686 => "01111101010111111111001100100110",
    687 => "11101111111001011010101010101100",
    688 => "11111010111111101111101100111011",
    689 => "01111101011011100001100101100100",
    690 => "11111111001111010110000010001111",
    691 => "01011100101101110111001101000111",
    692 => "11001110110111101010010000111001",
    693 => "11110111110111111001001110100100",
    694 => "01101101111111011001000001101011",
    695 => "00110011100000001011111001010110",
    696 => "00110110111001011000110110111001",
    697 => "11111110111111010101011100000010",
    698 => "00111111111111010011100001011001",
    699 => "00111111111000011101001101011011",
    700 => "01111110011101110101001111111010",
    701 => "01011111011111011011011101100101",
    702 => "10011111100011101100010001111011",
    703 => "00111111110100111011111111100110",
    704 => "01110101011111111011011111000101",
    705 => "01110101011101101111101000011000",
    706 => "10111111101111011101001100111110",
    707 => "01111011111111110000001111111101",
    708 => "11101111010111111101011011101100",
    709 => "11110111101010110110011100101010",
    710 => "11111101111111000101100010100010",
    711 => "11101111101101100001100110101001",
    712 => "01110010010101111011100101100001",
    713 => "11101100101111001100101001000001",
    714 => "00011110111111110111110110000011",
    715 => "01110100111110110000101011000011",
    716 => "01101111110110100110110101110000",
    717 => "00110011111011110000010110110001",
    718 => "11000111101110111110100101010000",
    719 => "10100111100101100110100110101101",
    720 => "01110011110101010010100110110111",
    721 => "10111101111111011111000110000001",
    722 => "11011101111011110110000010100000",
    723 => "11000111110011100111011111001001",
    724 => "11011101011011111010101101110110",
    725 => "11011101011111111011110010101110",
    726 => "01110111001111101000000000001111",
    727 => "01001110010100010001011100100010",
    728 => "10110100111111010000001011001100",
    729 => "01101101100100000110100010001011",
    730 => "11011111011111110101011101010010",
    731 => "01001001101110110000011111100110",
    732 => "01110111110100111001010011010111",
    733 => "10111111101110011101010101011000",
    734 => "11001110111110011011101110000100",
    735 => "00111111101101010100100010100110",
    736 => "11111110011011111000111101000111",
    737 => "00111011111111111110001111101111",
    738 => "11101111110111111001000011011010",
    739 => "00110001111010011111111111011101",
    740 => "01011110111111110001011010101101",
    741 => "00011001111110100101101100111001",
    742 => "11110011111101111010101110100101",
    743 => "01110101101100110010011100001010",
    744 => "10111001111011010100010001110001",
    745 => "11011111110111111011111011111111",
    746 => "10101011111110000001001100111000",
    747 => "11111010100110001001011111010111",
    748 => "01111100110100011010111101101010",
    749 => "00111110101110010110111110000000",
    750 => "01011011011011110011110011111111",
    751 => "01111101111111011111010000001100",
    752 => "00011011101111111101111011000011",
    753 => "01111011111111111001000001001011",
    754 => "01111011111110100010010000110100",
    755 => "01111011111111101111110111000001",
    756 => "10010111111101111011000100100011",
    757 => "11111101100101001100100110011010",
    758 => "10011111100110100011100100100110",
    759 => "01101100111111111100111011011101",
    760 => "01100111101101010010100101010010",
    761 => "01111101111111000011010011101111",
    762 => "11101100010111111011101000001111",
    763 => "00101001111111111101100111001100",
    764 => "01010110111010110010001100001011",
    765 => "10011100111110100111110011111110",
    766 => "01111011111010111110010010100101",
    767 => "11101011011111010001010111000110",
    768 => "11101111010111110111101111000101",
    769 => "10111111111111111111110101100110",
    770 => "11111011001101111110001000000010",
    771 => "10010011001101011110101100110111",
    772 => "10110110111101111001001010101000",
    773 => "11001011110011111000100010111001",
    774 => "01011101101111011011111001001010",
    775 => "10111111111001100011000101110111",
    776 => "01011110100010111010000111101001",
    777 => "00011111111010001011010010010001",
    778 => "11011011101111111111000011111100",
    779 => "00011111110000101000111111110011",
    780 => "01111011111111100101110010100000",
    781 => "01111010100011101010110011010011",
    782 => "11111110110101111010101110110001",
    783 => "10110110111011010101010100101101",
    784 => "11101111111111110010000111111010",
    785 => "11101011111111000100101110111001",
    786 => "10101001011001111011001110100101",
    787 => "11111011111110110000001001001010",
    788 => "11100101100111111110111111100011",
    789 => "10111011111111110001100011110000",
    790 => "01011010011011110011100011101111",
    791 => "11011111110110100101000110100011",
    792 => "01011110011111101001111011101001",
    793 => "10001111111001011111100111000000",
    794 => "11001111101101111001111101101011",
    795 => "11111100001010111001011010100111",
    796 => "01000011111110111001010101101011",
    797 => "01000001011111000101011000010001",
    798 => "10101111011111111101001001010000",
    799 => "11110100011011111101100000000100",
    800 => "01011111111110111001111011111111",
    801 => "11100011111011111010110011100011",
    802 => "11111101110101100001001010001101",
    803 => "00101111111111110110000111011110",
    804 => "10111111110011110101000010100011",
    805 => "11110110011111100111010111100101",
    806 => "01110101110011100111010110100110",
    807 => "01101111111111101010100001111010",
    808 => "01101111111011101010010010110100",
    809 => "00111111110110111111100100011010",
    810 => "11111110101101110100001111110001",
    811 => "11011110100011110111111011010110",
    812 => "01011101001011111100111110100010",
    813 => "10100111111011100100010101000010",
    814 => "11111000010111110100010101110010",
    815 => "11111111011100011100101101100100",
    816 => "01111000110001110001111100010001",
    817 => "00111011111111111000010110111010",
    818 => "11101111101110110001010100001101",
    819 => "11111011110011101000001001100110",
    820 => "11111100011011000000011111110110",
    821 => "11110100111101111110011111001111",
    822 => "10001101111010110110011101110011",
    823 => "01101010110111011111100001010111",
    824 => "00111100010111011100011111011110",
    825 => "01101111111111011110111100010010",
    826 => "10111111101111011101011001001011",
    827 => "01011011100011011001011111011100",
    828 => "11111101111011110110011001011011",
    829 => "01111011101111111111001111100100",
    830 => "00111110111101111100000110111111",
    831 => "01000111011111011010101000000111",
    832 => "10101011111111110010111100010010",
    833 => "10110101011111110010010011000101",
    834 => "00111111111110110111010010101111",
    835 => "01111110011111101010100110000101",
    836 => "00110001111111111101110100101100",
    837 => "10110000111001100111000110000101",
    838 => "01110011101110000001000111001100",
    839 => "11101110111101111111011110010101",
    840 => "11100101111111110000001110100101",
    841 => "11110111111010110110110010111111",
    842 => "01100001111111100000101001111111",
    843 => "01001111101110100111010111110111",
    844 => "10100101001010110010000010000010",
    845 => "01001111111011111111000011000001",
    846 => "01111111011110010101011010000011",
    847 => "01100011000011010111001000000011",
    848 => "01001111111011111100000111101111",
    849 => "11111110111110010001000100000001",
    850 => "11010010111011100010010010110011",
    851 => "00111111011111110101101111010001",
    852 => "01010111111001111110001100011110",
    853 => "01011110011110110001111010010110",
    854 => "00111010111110111110001011010111",
    855 => "00111111011111010001100111000101",
    856 => "00101101110011010111111000010100",
    857 => "11111101010011111010000011100111",
    858 => "11110111111111100111001101010110",
    859 => "01101100001111111001100100010101",
    860 => "11101111111110100000011010110001",
    861 => "01111101111101101100100110001001",
    862 => "11001111011111001110111110100001",
    863 => "00110010101111101100011111100100",
    864 => "11111101110101110011011001101001",
    865 => "11010011011110111000001100101000",
    866 => "01100111110001110010001100010110",
    867 => "01111011111111101110010110100000",
    868 => "11001001011101110110100010110010",
    869 => "11110010110011010110001111101000",
    870 => "10011111101100110011000000111110",
    871 => "11111011001001011010000111110001",
    872 => "00111101010101111000101000101101",
    873 => "00111011011101111001001010001111",
    874 => "11111111010000110111100101011111",
    875 => "01011011111111000001001011011011",
    876 => "00010011011111010001000111110101",
    877 => "11011101111111111100111001100001",
    878 => "00011110111111100000001100011110",
    879 => "11001111111011101100011001110000",
    880 => "11111011110111111001011100000101",
    881 => "01111110111001111110110010001101",
    882 => "01110101101111110010101100110011",
    883 => "10101111000111110100010100011101",
    884 => "01110110010111110000110011001000",
    885 => "10111110111110111111001101001100",
    886 => "11111001111101111100010000000000",
    887 => "00111111111010101010000010111011",
    888 => "10111011111101110111001100111000",
    889 => "10101101011011011000000001001000",
    890 => "11111101111101100101111100000111",
    891 => "01110111011111110101001101110100",
    892 => "01101111111001010000111011111110",
    893 => "01111010001100010110011100011110",
    894 => "11101111001110111000000101000100",
    895 => "11011111111110001100100101001100",
    896 => "11011111011111100000100101100110",
    897 => "11111100111110100011110110001010",
    898 => "10100100111111011000010011001101",
    899 => "01001001110111010111101000101011",
    900 => "00111010111011100101111011101000",
    901 => "11111111001000001000011000101101",
    902 => "00010110011111101100111001111101",
    903 => "11110100110011110101011101001110",
    904 => "10111110011101010101010100011111",
    905 => "10101110100110110011110111000000",
    906 => "11101011110011111001001100001100",
    907 => "11111110111011111010100100111011",
    908 => "01111111011111110010010011111011",
    909 => "11111111010011111010011001100110",
    910 => "10111111111011011111000111000111",
    911 => "00111111111110011100010001011011",
    912 => "01101111111111101010110001111110",
    913 => "01111011001110111001000111110110",
    914 => "00111101111101110100000110010000",
    915 => "01011111111111011110010101001100",
    916 => "00111110110110110001111010011001",
    917 => "01110011101110011001010010011100",
    918 => "11111110010111111111001011101111",
    919 => "11001111101110110001110001001100",
    920 => "10111111011110010100111110010011",
    921 => "11111110111011111011100110000110",
    922 => "11011110111011111010100110000100",
    923 => "01011111111011110010001101001110",
    924 => "01110111101111111100110011001001",
    925 => "11111001011111101111111110110111",
    926 => "11111110001101110100010001100111",
    927 => "11111000101111111101101001001101",
    928 => "01101111110000111101001011011111",
    929 => "01010111011111110000101111010110",
    930 => "11110111011001111000010001100110",
    931 => "10110111110101010010010001111100",
    932 => "11111001000110110010110110111100",
    933 => "01111101111110110001011010111001",
    934 => "01111111010101011000101101110101",
    935 => "11011111100010101110111101100110",
    936 => "10111010111011101110001001011110",
    937 => "10101011111100101101001111010111",
    938 => "11110111001111111000011101101110",
    939 => "01110101101111111101101111001101",
    940 => "01010010101101111110010101011011",
    941 => "10111111101010011000011110111001",
    942 => "01011011110110000100100101001110",
    943 => "01011101011011100010101111101011",
    944 => "11111110111100110110111100000111",
    945 => "11011011111001110100011001000110",
    946 => "01110111100110100101001101010010",
    947 => "01111110110011110100110010011100",
    948 => "11111000001100011001010010101101",
    949 => "10011101001100111001110100010000",
    950 => "10111111111111010010110100000000",
    951 => "10111101111011110000101101010001",
    952 => "11110111110111100111111000010111",
    953 => "10011010110101110000100010100101",
    954 => "11101111101101011100001010100010",
    955 => "01001111010111111101101011110110",
    956 => "00100100110001001010110110101001",
    957 => "11011001100111101010010011110100",
    958 => "00010111111111110111100101101000",
    959 => "10111111111011101000100111100110",
    960 => "11011111001110101010011101111111",
    961 => "11110111000110110011001110110000",
    962 => "11111100110111010100011101000011",
    963 => "11100101111111011100110000101100",
    964 => "01111001111101110110001111000011",
    965 => "01101111110111100000011000110111",
    966 => "11100101010011110010110111011111",
    967 => "00110111100001010101011000110011",
    968 => "00011100110111010000111010100001",
    969 => "11101101110111110010010010000100",
    970 => "11110011111111110110001100110001",
    971 => "00111010001001100000110111011100",
    972 => "11011111010111011010101111000010",
    973 => "01110111111110010001110000100010",
    974 => "11000011111001110100011011110011",
    975 => "01111010111110110001001011100001",
    976 => "01011110111111111011011110111101",
    977 => "11000011111110110100001100000001",
    978 => "11101111111111110011111001111000",
    979 => "11100010101111110000001100101111",
    980 => "01011111111001110000100011100011",
    981 => "01110110110110110001000101010000",
    982 => "10111100011101110110110101000110",
    983 => "11110011110110111000000001011000",
    984 => "11100111111111111000010111101101",
    985 => "11110111111111110110001111111000",
    986 => "00001111111110101110101110110000",
    987 => "01110111111111110001101100001101",
    988 => "01111010000110110100010101100010",
    989 => "01011010010111111100101101110011",
    990 => "10011011001110101101110010100100",
    991 => "00111111101111011011001001101000",
    992 => "11111010111101010000011100011010",
    993 => "00001011010111111010111100010111",
    994 => "10111111111111101001001100011100",
    995 => "11100100011111010001001110110000",
    996 => "10101101111011011110111010111100",
    997 => "01011110001110100000101111101111",
    998 => "10101100010111110011110110111010",
    999 => "11110011111001111110110111001100");

  constant ans_lut : lut := (
    0 => "11101111111101010111011101101110",
    1 => "11011111011111011011001010010100",
    2 => "11011101101111111001011101101001",
    3 => "01111101111101111101011111110011",
    4 => "01101110101111111011100101011101",
    5 => "10101010101111110011010111011000",
    6 => "10010011101110110001110111110101",
    7 => "11001100111101100011010011001000",
    8 => "01111101010111111010011100000000",
    9 => "01111011011111110100111010110111",
    10 => "01111011110111010010111000111000",
    11 => "01101111100111111111111111011011",
    12 => "10110111100111110100111001001010",
    13 => "01011011011111010111010001111111",
    14 => "01110111111111110001101111001010",
    15 => "01011111101110110101000010100010",
    16 => "10010111001111100011011010000110",
    17 => "01101101111111111110110101010101",
    18 => "01000111010111100101100011010011",
    19 => "11010110101110101000011101110000",
    20 => "01011101011110110011110001100001",
    21 => "11110111001010011101000011101010",
    22 => "11110111111111110000111001001100",
    23 => "11111101100101110000010110000011",
    24 => "11110111111110110101000010011100",
    25 => "00011111111011111101100011010001",
    26 => "11101101110110011000011000000101",
    27 => "00110101110101100111101001100011",
    28 => "01001011111101010001010000110101",
    29 => "11101011101111110011010100001001",
    30 => "10111011011111101100111000111100",
    31 => "10100111011111110001100010101010",
    32 => "01111000101110111110011110100110",
    33 => "01111111010110110011100101000000",
    34 => "11110101111011010101110101100010",
    35 => "11101110011011100101010001100100",
    36 => "11101011101100111110011011001010",
    37 => "10101101010110111011111110110011",
    38 => "11011111110011110010000000001001",
    39 => "01111100110111100110110000111011",
    40 => "01111110111011111010111100110110",
    41 => "11101111111111110100011000101010",
    42 => "01101111001111111111010010011111",
    43 => "01011110110110111010010100011010",
    44 => "01111101110111101110101101111000",
    45 => "01110011010111111110100111101010",
    46 => "10101011101010110101110111011110",
    47 => "00110111101011111001100011001011",
    48 => "00001111110000110001100100111101",
    49 => "01111000111110110110101111100011",
    50 => "01101011111111001001100100001110",
    51 => "11010111110110111110100101000000",
    52 => "00011111011101101000010011000110",
    53 => "01011110111110111111011110001011",
    54 => "01001011111111111100001000010000",
    55 => "01111110101111110010010101010000",
    56 => "01011011011010110101010010110110",
    57 => "11000110111111100111100110001010",
    58 => "11101111111111011000100000101111",
    59 => "01100111011011110001001101001100",
    60 => "11111101111101011000011010011111",
    61 => "10011111111011101010000101001110",
    62 => "00111011111110110010110000000001",
    63 => "11110111111111111001111100000000",
    64 => "11011010111001000001101010011110",
    65 => "01110011101111000001111000110000",
    66 => "11100111011100111001011011010000",
    67 => "11011111100111111011100011110110",
    68 => "01110010111010111001111111100111",
    69 => "11101011111111111110011010001000",
    70 => "10111111110110100011110000011101",
    71 => "01111011110110110001100010100110",
    72 => "00110110101111111101011001000011",
    73 => "11011111011101111101000100000001",
    74 => "01111101010111111111010110100100",
    75 => "11111101010111110100010010000001",
    76 => "01101101110011110101100111000010",
    77 => "00111111111010111001101110101110",
    78 => "10111110111111110111000010101010",
    79 => "00001011111110001100101100000010",
    80 => "01111011001101100100010110010010",
    81 => "01011110011100110011111011110101",
    82 => "01111100110011111111011111111010",
    83 => "01011111100111101010100001101101",
    84 => "01100100110010111111001010000001",
    85 => "11001011001111111110101001011010",
    86 => "01000110110111100111010101011110",
    87 => "11100111011111111001110101010111",
    88 => "00111010111111110001111100010001",
    89 => "11101111110111110010101010101101",
    90 => "01010110011111110000111100111111",
    91 => "00101010111111010100100101100001",
    92 => "01111011100111000000101000110010",
    93 => "11111011111011110100010101010100",
    94 => "01100100010110011011111001100111",
    95 => "00101111001111100000011110010001",
    96 => "10100101111110110011111110010100",
    97 => "11111010011101011101111000001101",
    98 => "01101110111101110000100100101100",
    99 => "01011111111100111000100100000101",
    100 => "00111101101111111100010011101010",
    101 => "11111101110111110000101110101000",
    102 => "11110111000011110111010000000110",
    103 => "11111110011111100010011110111011",
    104 => "10101111011111110000111100010110",
    105 => "11111110111010100101001101101101",
    106 => "11011001110101010011100010000100",
    107 => "11100101001101111101100010110100",
    108 => "11110100111111111100000011011111",
    109 => "11100010011111000011111110100000",
    110 => "11011101111111110111100110001011",
    111 => "01111110111101110011001010001001",
    112 => "01001111101111100100101001011001",
    113 => "11111110111111011011010111000011",
    114 => "11011101011101110111011111100011",
    115 => "00100110111110111010100000000001",
    116 => "01111011011111110110100111001000",
    117 => "00100011110011111101101101100100",
    118 => "01111100000111100000110101000100",
    119 => "01011111011011111110001001100010",
    120 => "10100011101011110000100100000001",
    121 => "01110011101011101100111010010111",
    122 => "10000011011110110011111110110000",
    123 => "10110101111001010000010101000011",
    124 => "10000110100001110111000011100111",
    125 => "00111011110100111001010011011111",
    126 => "00111111110100001100110010110001",
    127 => "00000111111101110111001100101001",
    128 => "01101111111111111100111011101010",
    129 => "11011111111111011010110000111101",
    130 => "11010111001111110000010001010001",
    131 => "11111110011110011100110111000111",
    132 => "00111011111110110100111110101110",
    133 => "11111110111111110001000001100101",
    134 => "01110011111001110101110101000011",
    135 => "11111111011111000010101100010101",
    136 => "11010110111110111110100011010000",
    137 => "01101110101100111111101011001110",
    138 => "11101011101101010111101000111111",
    139 => "10111111100111111111010010011001",
    140 => "01010001010111100010011011110101",
    141 => "00111011001111101011101100101111",
    142 => "00111110100110110100001110111111",
    143 => "01101111111111100100000111111110",
    144 => "11100111011011111101000011100110",
    145 => "00011110101011010100010000111011",
    146 => "00111011111110011011010001101000",
    147 => "01010100110111110100011111011000",
    148 => "00110111110110111111000011011011",
    149 => "11011011111101011011011110010101",
    150 => "01011100010111110000101101011111",
    151 => "01111110001011110001010110011110",
    152 => "10111010011011110010000011011001",
    153 => "00011011101110101110001001000011",
    154 => "01110111111111100111110000100001",
    155 => "00100011011101111010101000110110",
    156 => "11100111111011111001100000100110",
    157 => "01011111111011110011110100110101",
    158 => "11111111001101111110111101111110",
    159 => "01001111011011011100101111100010",
    160 => "10110011100111111100010110000010",
    161 => "00111110111011111010010000000111",
    162 => "01111100111001110011111010110111",
    163 => "01110111110111110100110000000110",
    164 => "01101111111101111100001010101011",
    165 => "01101111111101010100101110010101",
    166 => "10101101111110001101011011011101",
    167 => "11111110111111110111111010011100",
    168 => "10111000110110110000010010110100",
    169 => "00111101110110111111011000010101",
    170 => "11010110111110101011001001111101",
    171 => "11110111111111110011111000011100",
    172 => "00111111111111110101010011000000",
    173 => "01111010111111111111000111101001",
    174 => "10110111111111110100010000011001",
    175 => "00110111111111101000110110101001",
    176 => "10111110011111110010011011101101",
    177 => "01101111101110111110011110000110",
    178 => "11111111010110110000010011101110",
    179 => "01011011110011001100110100011101",
    180 => "11001111111110010110000011110100",
    181 => "11101101101011110010111011001010",
    182 => "11101110111111110111010010001100",
    183 => "10001010101001101000000001111100",
    184 => "01111110111111011011111111100110",
    185 => "11011111111101111000001010100101",
    186 => "11110101110011110101101111000110",
    187 => "01011111111101100000110101101101",
    188 => "00011011100111111010010100101111",
    189 => "01101100101111010011000000000000",
    190 => "11010111111011101101100110010100",
    191 => "01111110110110101011010110110100",
    192 => "00011011111110110100101010100001",
    193 => "00101011111101111011101001001110",
    194 => "01111101011110111100111010001011",
    195 => "11011111011111110001000100111110",
    196 => "10111011110100110000110111111000",
    197 => "11111111011101100100010111011100",
    198 => "01010111110110101000111100000101",
    199 => "11101110111011110111000011001000",
    200 => "01111011111011111000010011110000",
    201 => "01100101111101110110001110010010",
    202 => "11111111001010111000000010010111",
    203 => "00110111110101110000110000010111",
    204 => "01110111111110111101100101000111",
    205 => "01101110111111111100100000011101",
    206 => "10111011111111101100010000101101",
    207 => "01111111011111011011111001010100",
    208 => "01011111101101110110011110010101",
    209 => "11110101100111110010001101110000",
    210 => "11111111010111001110001101010011",
    211 => "11110011111111111101101110101111",
    212 => "11011110111110000010111110100101",
    213 => "01111110100101111100000101000101",
    214 => "11101110110111110011111111100110",
    215 => "00101111111111101001010101001100",
    216 => "11011111111110111001010111010111",
    217 => "00101011111111101011010100001110",
    218 => "00111110110101111100011001111010",
    219 => "11001111111101110001110101010001",
    220 => "10111111001111111010000101010110",
    221 => "10111111110111010000111101110111",
    222 => "10110111111001110010111100111100",
    223 => "11010011100011111010011101100101",
    224 => "01011011011101011001110000110100",
    225 => "11110111011111011100111110001101",
    226 => "11001111011101111000000001101110",
    227 => "10111111111110110110101100000101",
    228 => "11110111110111111011011101010101",
    229 => "01111011011111111010001011001011",
    230 => "11101010111111001111101010111001",
    231 => "10011111101010111000000010110000",
    232 => "10111011101001100111011000101011",
    233 => "11010011111111110100011100101001",
    234 => "11110111101100011000000110110000",
    235 => "01111110111011110111001001000110",
    236 => "10011001111011101000100110001000",
    237 => "10110111111111011100001101111100",
    238 => "11111110111001011001110011000001",
    239 => "11111101111111111111000110010101",
    240 => "11110110000111101000111010010010",
    241 => "01111001111101110111101111000001",
    242 => "10110111100111111000011110111111",
    243 => "00111111010111011111101001110011",
    244 => "01011111011111101001111101111010",
    245 => "00011010101101111010010101110110",
    246 => "10110111011101111100011110100011",
    247 => "01111001011101110100100000101101",
    248 => "01011001111111100111111000111101",
    249 => "01111110101101110101000000001000",
    250 => "01111001111101110111101011001010",
    251 => "10111111010111110000101000101111",
    252 => "00111110111101011111111101001101",
    253 => "01111001111111111000011010101011",
    254 => "10011111001111110001001100111110",
    255 => "00001110111111110110001011100110",
    256 => "01101111101001010000111011010100",
    257 => "11101011111001111100001000010110",
    258 => "11101101110110101001111000000011",
    259 => "11011111111110111010011010000110",
    260 => "11101110011110011111101111000011",
    261 => "01101110110010010110100110100000",
    262 => "01111101110111101010101111110111",
    263 => "10101110011101101010011101100111",
    264 => "01110111011011110111101110101100",
    265 => "01111110111111110001101010111000",
    266 => "10110101111111111101000100000000",
    267 => "01010101010111110011010010111101",
    268 => "01011111001111111100000100101111",
    269 => "11101110101101101101000010100101",
    270 => "10111011111111000000111010111011",
    271 => "01111100101111101110100011000000",
    272 => "00101111110101111001000110111100",
    273 => "01111101011111111111000000111000",
    274 => "01101110111111110000101110100110",
    275 => "01111111010111101101001110011011",
    276 => "01101011110111110111110111001001",
    277 => "01111110100111100001001100111011",
    278 => "01011111001110110111101110100011",
    279 => "10111110111110111011111000101001",
    280 => "10111110111111110101110001101011",
    281 => "01101111001001110001110001100011",
    282 => "11101101111111111001011000010011",
    283 => "00111011101110100111101110100110",
    284 => "00110111011011100110011001110011",
    285 => "11110111000111100011110011101001",
    286 => "10010100100101011001101000001101",
    287 => "11110100011000111111100101101100",
    288 => "11110111111111111111111011011000",
    289 => "11110011001110110001111110111010",
    290 => "01011111111111010010100110111011",
    291 => "00010111111110111111000100100110",
    292 => "01101111111110011101100000110000",
    293 => "11111011010110011101011000111100",
    294 => "01111100110110101101101110001111",
    295 => "10111111111110111010100010111110",
    296 => "01101101001111011111101100010101",
    297 => "01111101111111110010011000100010",
    298 => "00111011111111011101000110111100",
    299 => "11111010011011110010010010101010",
    300 => "11111001100111010101100011101111",
    301 => "01111011111111101010101001001001",
    302 => "00100111111111110111001000011001",
    303 => "00001111100111110001101011101011",
    304 => "11111110111011111000001100000101",
    305 => "11111110011010110010001001110111",
    306 => "01111110111001111101110001010000",
    307 => "01111011110011010010001101111011",
    308 => "01111111011110110011001111000001",
    309 => "00101111111011110011011100000110",
    310 => "11011101001110001010000110100000",
    311 => "11111011110111000011001100010010",
    312 => "11010111101111111111111011110001",
    313 => "11010111111101001010101110001011",
    314 => "11010111110111011011100101010001",
    315 => "11101011011010100100101011011100",
    316 => "01111010011111001111100110001011",
    317 => "10110110011111101001110001011011",
    318 => "10111111011001100011100101010101",
    319 => "11111011111111100101100100011101",
    320 => "10111101011011111001001110001100",
    321 => "00011011011101111110011111111011",
    322 => "00111110111100001011011000010010",
    323 => "01101111100111110110011010110100",
    324 => "10101001011111100011000010111011",
    325 => "11100111111011110100101001000001",
    326 => "11001111001111110111101110110000",
    327 => "11110111001111111011101110001010",
    328 => "11110111111110111010000100010011",
    329 => "01111011111011110111110100010000",
    330 => "11110110101111111010000001000101",
    331 => "10111100101101111001111000101011",
    332 => "01011111101010011000101100010010",
    333 => "01101111101111110101110000000001",
    334 => "01101111101011110011001101001101",
    335 => "11011101111111111010011010010101",
    336 => "11111110111001110001001111110110",
    337 => "11111011111110101001000001101001",
    338 => "01000101011111100100100111000000",
    339 => "01011101100101011000001011111110",
    340 => "01111110101011110010010011110001",
    341 => "01110110111111101101110100110011",
    342 => "11111110111001110010010111101010",
    343 => "01110111111110110101010101010111",
    344 => "01110101101111110110101000110110",
    345 => "11001010111101010001100110010110",
    346 => "01110110101110110011001000111110",
    347 => "00011110011111111101111111100010",
    348 => "11011011011101101000100011010111",
    349 => "01101110011101010111110111001101",
    350 => "01110011111010011010010000001101",
    351 => "11110100111101111000000100001001",
    352 => "01011011111011010010101110010010",
    353 => "00111110111100011111010110011010",
    354 => "11011110111011000101111011001010",
    355 => "01011111001110111111101100001000",
    356 => "11011010110111111011101001000100",
    357 => "11101100111110100111011000100100",
    358 => "01101111101111100100010111111100",
    359 => "11111000001111110010110011011100",
    360 => "10011110111111100011010001100010",
    361 => "01111110011101110001111111101110",
    362 => "01111100111110110101111110101110",
    363 => "11100111111111111010100010101001",
    364 => "11101011101110110110110111001000",
    365 => "01111011011110110011100000110010",
    366 => "11110011110011110100011111101011",
    367 => "01110111001111110100100001011001",
    368 => "11110011111000011000111101000100",
    369 => "11001001111111111100100001010100",
    370 => "10111110011111111001001111000000",
    371 => "01111001101111110110111000000011",
    372 => "00111111111111111100111000110010",
    373 => "11100111100111110101000111110111",
    374 => "11011110011111111010011110011110",
    375 => "10011111011111101101110010111000",
    376 => "01010111011001111000010001101100",
    377 => "01110010111101010010001100111000",
    378 => "11011111111110111010111100010100",
    379 => "01100011110110101000101110001111",
    380 => "01010011011110101000100100111000",
    381 => "01010111100101011111011011010110",
    382 => "01110111011110111100100010100101",
    383 => "00110000111110110001010011110010",
    384 => "00101001101110101100111110100100",
    385 => "00111101111101111000001001101111",
    386 => "01010101011101111101100010000111",
    387 => "01101100001001011010000000111001",
    388 => "11101111001111110010110011011000",
    389 => "10001001101101010100011110110001",
    390 => "01111100000111100111111110000100",
    391 => "01101111111111111000111011110010",
    392 => "10111110100011101011111001010010",
    393 => "00011111111111111110000110010110",
    394 => "01011011111011010001110101011100",
    395 => "01100110010000010101100011110000",
    396 => "10101111111011000111011011111011",
    397 => "11110111111011110001011010010101",
    398 => "00011011100101000110101111010011",
    399 => "11011111010110111110010000010011",
    400 => "00000110010011110110110101101011",
    401 => "01111110011001001100010001111111",
    402 => "10111100111110011110010001010100",
    403 => "11110011110111101010001111010101",
    404 => "11111010110101111101100001001111",
    405 => "01010111111111010000011010010100",
    406 => "11101101101111010111000011001110",
    407 => "11111111011111001110000010000011",
    408 => "01111101000111110010101011010001",
    409 => "01001011111110011110001111100000",
    410 => "11101011100010111011011110000101",
    411 => "11101011111110111010000101001010",
    412 => "00001101110111010000001010001000",
    413 => "11111101001100110000100110101001",
    414 => "01101111111111110000101000110111",
    415 => "01101111101011100011100001100100",
    416 => "10011111101110110101000111010101",
    417 => "11011010111111101110000011010100",
    418 => "11110101111000101010011101010100",
    419 => "00011111111101110101110100100110",
    420 => "01111001110100011010010000000110",
    421 => "01111110110110011000010110110110",
    422 => "11111001101101111100111001001101",
    423 => "10100111011111000101100000110001",
    424 => "10011111111101111100010001110011",
    425 => "11100101111111111000101010111111",
    426 => "00011101010001110011001100010000",
    427 => "01011110110101111110101100011010",
    428 => "01110100110001111111110100111011",
    429 => "11001111111100111100011011110110",
    430 => "01111111010110101110001011000001",
    431 => "11110101100111111011010101111111",
    432 => "00110111110111110001000000001101",
    433 => "01110111011000111000110100000000",
    434 => "01101110001011101110011111110101",
    435 => "01001111111111110011111100111001",
    436 => "01010111111101101101001101101000",
    437 => "00100001111111010101101011010011",
    438 => "00110011110111110010111010000111",
    439 => "01110110111110101100001011110001",
    440 => "11011111101110111100001010111100",
    441 => "01111101110011100101100010110111",
    442 => "11110111110100111101101011111000",
    443 => "01111100011100111001000010001111",
    444 => "11011111111111110011100010010100",
    445 => "00010111011101010101011011100000",
    446 => "11100110111011100100111111101100",
    447 => "01011110111111010010101101111000",
    448 => "11010111111111110001111001010000",
    449 => "11011111111010111100011100010011",
    450 => "01111011011111111001111101101000",
    451 => "01111110011111100010001001111001",
    452 => "11010011000110000011110000110000",
    453 => "01111111001110111010110101000001",
    454 => "01111100101110010100110011010011",
    455 => "10111111111111110110010111001001",
    456 => "01110111010111011110000010000010",
    457 => "10011001110101111111111111111111",
    458 => "01011111111001110100110111011110",
    459 => "00100100111111110011010001101100",
    460 => "01010100111110010111010011001010",
    461 => "01111101010110100000101110101101",
    462 => "11101110010110101011001110101111",
    463 => "11010111110111111000011110000110",
    464 => "00111011000001011100001011010011",
    465 => "10111111111110111111111000100101",
    466 => "11101011111111110110101010010001",
    467 => "01111011010110111101101110101100",
    468 => "00111110111111110111001011000100",
    469 => "11110010110100111100011010110011",
    470 => "10011100100110011101010101000110",
    471 => "11001011111101110101001001101000",
    472 => "01100111111110111011100101010000",
    473 => "01010101111111011000111000001011",
    474 => "01101111111111010110011101110100",
    475 => "11111111011100111110111011111010",
    476 => "11110111101001110001011110101000",
    477 => "01011111011111110110111000111010",
    478 => "10111111110010111101100101111110",
    479 => "01010111111011011011011000100010",
    480 => "11110110111101010101101001111100",
    481 => "10111111101011110010001010011100",
    482 => "01010111111000111111000100001110",
    483 => "00110111110000111111001001011000",
    484 => "01011111111111110000100000100011",
    485 => "11011110110010111100110001010011",
    486 => "01101101111111111101000101010000",
    487 => "11111111011110110010000110111101",
    488 => "01011111011110110100101010100001",
    489 => "10111111100110110100111010101011",
    490 => "11110110111110111010010001010100",
    491 => "10010010101011111011000000011100",
    492 => "01111100111111110100000011001110",
    493 => "10111111010111011100111000011101",
    494 => "00000100111111111110110000011111",
    495 => "11000111110111111111000111110001",
    496 => "10011111101011111010010011110011",
    497 => "00011111100101100111110011000100",
    498 => "11101111001111111010100111101110",
    499 => "00110011100110010100110111000011",
    500 => "10011011101101110011011010111010",
    501 => "10001010011110110000110010011101",
    502 => "11111110010110101001111110111010",
    503 => "01111010010110110110011101100110",
    504 => "00110110011111101011011110001100",
    505 => "11011011111100010010001111110110",
    506 => "01011101110111110001110001100101",
    507 => "11111101001101110110111001101111",
    508 => "10111110110111011010010010110000",
    509 => "01110000110011110111011110000001",
    510 => "11101111111111111101011101101011",
    511 => "11010101111011110111110111111111",
    512 => "11011111100001111100001101001100",
    513 => "01110111100111100110001110011011",
    514 => "11010111111111110000001000010001",
    515 => "11111001111111010001010011110110",
    516 => "01001110101010101110110110110000",
    517 => "11010101101011110001111110001010",
    518 => "00110111111110111110010110111010",
    519 => "00111110011110101001100100100011",
    520 => "11110110111111101101001101011111",
    521 => "01010101001111110001101100111010",
    522 => "01111011101001010111101000010110",
    523 => "01111001010111111111100111101010",
    524 => "01110101111111010100011011010100",
    525 => "11011011001100110010000000000011",
    526 => "01111010010110110011111100110001",
    527 => "01111010111111000000010000100111",
    528 => "11000110111111011110000010011110",
    529 => "01111101100111111010011000100010",
    530 => "01011111110111100110111110110000",
    531 => "01011111111111101100001000010111",
    532 => "01111110011111111010010101111001",
    533 => "01101011001101111100101100101010",
    534 => "11101101010011011000000101001101",
    535 => "11010110101011110001010110011110",
    536 => "10111001110111010111010011110010",
    537 => "01111111011010001110100011010111",
    538 => "01100011111011010010001101111101",
    539 => "11101111011100111110011100011110",
    540 => "10110111111000101101100001101101",
    541 => "10010111111111110111010001110010",
    542 => "11111011100111110000000100100100",
    543 => "01111011110100111011101001101011",
    544 => "11101100110011010111111011010001",
    545 => "01111110100101101101011101011000",
    546 => "00011111011111111111010001011111",
    547 => "01011101110110110111110110111100",
    548 => "11001101111011111000001111101010",
    549 => "10000111001101110010010100001100",
    550 => "11111011111110111010110100110100",
    551 => "10111110111001110101100111100011",
    552 => "11000110101111100110101110000010",
    553 => "01011110111111110001000100101110",
    554 => "01111101010011010010010101111011",
    555 => "11111101111011111111111101101111",
    556 => "10101010111101110001010110000111",
    557 => "01001111111101101110011001011100",
    558 => "11100111001011011110001001010110",
    559 => "01111101101011100011000001111111",
    560 => "10100110110111110101001110101111",
    561 => "01110001011111100101001100011110",
    562 => "01110111000011111011111010111000",
    563 => "01100011110111000001101001010010",
    564 => "01010111101011111101110000111111",
    565 => "11111110001101110001111001101111",
    566 => "01101101111110011110100110101100",
    567 => "01111010111110110111100011011100",
    568 => "01111110111111110001100011110001",
    569 => "11011111011101101111001100101000",
    570 => "01110111101111111001110001000000",
    571 => "00111001110110111000000000000101",
    572 => "11101110111111011111001100101010",
    573 => "01110111100010111000000110111010",
    574 => "00110011011110111100101110001110",
    575 => "10011111101111111000111100101111",
    576 => "01110111010111111101011100011001",
    577 => "01111101111110011111000010101010",
    578 => "11101010111111111011100101010101",
    579 => "01011111111111110111100110010101",
    580 => "00011000111001111101001010000011",
    581 => "01111111011111111100101110110110",
    582 => "11100111111100100010000111110110",
    583 => "10111011111011111011011100001010",
    584 => "01101111001101101110001011101010",
    585 => "01011101011011101001110011001001",
    586 => "01101111111111000011000011110010",
    587 => "00110011111111010011001110001111",
    588 => "01111111010111010110010101110101",
    589 => "01110110101001110110010011100111",
    590 => "10111110110011100001111001011011",
    591 => "10001111111101011101011011110010",
    592 => "00110110111001111101000111010001",
    593 => "11101011011111100001101000000010",
    594 => "01111100111001110010010111011100",
    595 => "01110101111100101110001101101011",
    596 => "10011101111110111010100010110100",
    597 => "11011111101111110011011000100101",
    598 => "11011011011011110100000001001000",
    599 => "01011111111101110000100111110001",
    600 => "00101110111111111001100000111001",
    601 => "01011101101111110101101010011111",
    602 => "00001111011111110011011010101111",
    603 => "00011111011111010111101111011001",
    604 => "01100011110001011000110101001011",
    605 => "00101011101101111001000011001000",
    606 => "01101111100110111011101010101100",
    607 => "01111101101111101111100000000010",
    608 => "11011111111111100011100111110111",
    609 => "10011111011100111100000100110011",
    610 => "11101001111010100000111101110000",
    611 => "11000111111111010010001011000011",
    612 => "11110011111110111100100110100111",
    613 => "01111011100111010101111010100100",
    614 => "01111110110111101111000001111100",
    615 => "00110111011100101100000000001010",
    616 => "10111111111001111101100101001001",
    617 => "11101111100111010100110100100110",
    618 => "11111101011111110001001000111100",
    619 => "01101100111111100100010110101001",
    620 => "10111101101110110010011111110100",
    621 => "11100111111110111010000110010111",
    622 => "11111010110110110101101110001001",
    623 => "11101010111110110111111101001110",
    624 => "00101110100100111100110010110010",
    625 => "00010111110110011011000010001111",
    626 => "10001111001101010000010100011101",
    627 => "01100100111101110000011000010010",
    628 => "01111110110111100100000010110101",
    629 => "11111011111111111001010101001000",
    630 => "01110010111111100000000111111111",
    631 => "11111110101000111000000010010011",
    632 => "00110011111111111100000001011101",
    633 => "10011110100011110101100000000101",
    634 => "11011011010111110100001110110010",
    635 => "00011111001111111110000111100100",
    636 => "11101001101100100110010000011001",
    637 => "11110100111011100000101000110110",
    638 => "01111011111001110000001101000100",
    639 => "11111100111010111100011100100101",
    640 => "11111001111101111100100111111001",
    641 => "01010101111111111111110111111010",
    642 => "11111110101111110001010101011101",
    643 => "00111011101111111001011000100111",
    644 => "00011010011001100101100010101110",
    645 => "01011111010010011000110100010011",
    646 => "11101111110011010110110000010001",
    647 => "01001011111011110101001101111000",
    648 => "00111111011011111000111011000110",
    649 => "11111001101110111100110100011000",
    650 => "11111111001101010011011001100110",
    651 => "11101001110111001101000111011101",
    652 => "01010111111010110110000111111101",
    653 => "10111101001110111111101101100010",
    654 => "01100111010111111101110110000010",
    655 => "10101111111011100001101000101100",
    656 => "11111010110110100001101000111100",
    657 => "00111111010111001100001110110101",
    658 => "01111010011011011111010011000001",
    659 => "11111010011111011000100101001011",
    660 => "10011010110110011000001111110110",
    661 => "11110111101111101101111101100011",
    662 => "11011101110011101000100010111100",
    663 => "11011111110110101000001000111111",
    664 => "01101100111111010101011001100110",
    665 => "11110101110011010010111110111011",
    666 => "10001101011111110000110101100000",
    667 => "11101111111110100001011100100100",
    668 => "01111100100011111110100010111011",
    669 => "10101111111101111101011100110010",
    670 => "01110001111111101101100000011001",
    671 => "00011111111011110111010111000010",
    672 => "01011001110111101001100010111110",
    673 => "01011101111111110001011001001100",
    674 => "00111111100111110111101000001011",
    675 => "01111110011111011101010110111000",
    676 => "00111111001111011011011110101000",
    677 => "11000110011011010100111100001111",
    678 => "01011101010111101100101011100110",
    679 => "11100101111111111001101011111111",
    680 => "01011010111111111011010110001011",
    681 => "01011010111010110111001100010101",
    682 => "00011111101110011101011111111000",
    683 => "01001000101111110010101010000110",
    684 => "11001011101110100011011011000100",
    685 => "11011110111111011100001110011011",
    686 => "11111101010111111111001100100110",
    687 => "01101111111001011010101010101100",
    688 => "01111010111111101111101100111011",
    689 => "11111101011011100001100101100100",
    690 => "01111111001111010110000010001111",
    691 => "11011100101101110111001101000111",
    692 => "01001110110111101010010000111001",
    693 => "01110111110111111001001110100100",
    694 => "11101101111111011001000001101011",
    695 => "10110011100000001011111001010110",
    696 => "10110110111001011000110110111001",
    697 => "01111110111111010101011100000010",
    698 => "10111111111111010011100001011001",
    699 => "10111111111000011101001101011011",
    700 => "11111110011101110101001111111010",
    701 => "11011111011111011011011101100101",
    702 => "00011111100011101100010001111011",
    703 => "10111111110100111011111111100110",
    704 => "11110101011111111011011111000101",
    705 => "11110101011101101111101000011000",
    706 => "00111111101111011101001100111110",
    707 => "11111011111111110000001111111101",
    708 => "01101111010111111101011011101100",
    709 => "01110111101010110110011100101010",
    710 => "01111101111111000101100010100010",
    711 => "01101111101101100001100110101001",
    712 => "11110010010101111011100101100001",
    713 => "01101100101111001100101001000001",
    714 => "10011110111111110111110110000011",
    715 => "11110100111110110000101011000011",
    716 => "11101111110110100110110101110000",
    717 => "10110011111011110000010110110001",
    718 => "01000111101110111110100101010000",
    719 => "00100111100101100110100110101101",
    720 => "11110011110101010010100110110111",
    721 => "00111101111111011111000110000001",
    722 => "01011101111011110110000010100000",
    723 => "01000111110011100111011111001001",
    724 => "01011101011011111010101101110110",
    725 => "01011101011111111011110010101110",
    726 => "11110111001111101000000000001111",
    727 => "11001110010100010001011100100010",
    728 => "00110100111111010000001011001100",
    729 => "11101101100100000110100010001011",
    730 => "01011111011111110101011101010010",
    731 => "11001001101110110000011111100110",
    732 => "11110111110100111001010011010111",
    733 => "00111111101110011101010101011000",
    734 => "01001110111110011011101110000100",
    735 => "10111111101101010100100010100110",
    736 => "01111110011011111000111101000111",
    737 => "10111011111111111110001111101111",
    738 => "01101111110111111001000011011010",
    739 => "10110001111010011111111111011101",
    740 => "11011110111111110001011010101101",
    741 => "10011001111110100101101100111001",
    742 => "01110011111101111010101110100101",
    743 => "11110101101100110010011100001010",
    744 => "00111001111011010100010001110001",
    745 => "01011111110111111011111011111111",
    746 => "00101011111110000001001100111000",
    747 => "01111010100110001001011111010111",
    748 => "11111100110100011010111101101010",
    749 => "10111110101110010110111110000000",
    750 => "11011011011011110011110011111111",
    751 => "11111101111111011111010000001100",
    752 => "10011011101111111101111011000011",
    753 => "11111011111111111001000001001011",
    754 => "11111011111110100010010000110100",
    755 => "11111011111111101111110111000001",
    756 => "00010111111101111011000100100011",
    757 => "01111101100101001100100110011010",
    758 => "00011111100110100011100100100110",
    759 => "11101100111111111100111011011101",
    760 => "11100111101101010010100101010010",
    761 => "11111101111111000011010011101111",
    762 => "01101100010111111011101000001111",
    763 => "10101001111111111101100111001100",
    764 => "11010110111010110010001100001011",
    765 => "00011100111110100111110011111110",
    766 => "11111011111010111110010010100101",
    767 => "01101011011111010001010111000110",
    768 => "01101111010111110111101111000101",
    769 => "00111111111111111111110101100110",
    770 => "01111011001101111110001000000010",
    771 => "00010011001101011110101100110111",
    772 => "00110110111101111001001010101000",
    773 => "01001011110011111000100010111001",
    774 => "11011101101111011011111001001010",
    775 => "00111111111001100011000101110111",
    776 => "11011110100010111010000111101001",
    777 => "10011111111010001011010010010001",
    778 => "01011011101111111111000011111100",
    779 => "10011111110000101000111111110011",
    780 => "11111011111111100101110010100000",
    781 => "11111010100011101010110011010011",
    782 => "01111110110101111010101110110001",
    783 => "00110110111011010101010100101101",
    784 => "01101111111111110010000111111010",
    785 => "01101011111111000100101110111001",
    786 => "00101001011001111011001110100101",
    787 => "01111011111110110000001001001010",
    788 => "01100101100111111110111111100011",
    789 => "00111011111111110001100011110000",
    790 => "11011010011011110011100011101111",
    791 => "01011111110110100101000110100011",
    792 => "11011110011111101001111011101001",
    793 => "00001111111001011111100111000000",
    794 => "01001111101101111001111101101011",
    795 => "01111100001010111001011010100111",
    796 => "11000011111110111001010101101011",
    797 => "11000001011111000101011000010001",
    798 => "00101111011111111101001001010000",
    799 => "01110100011011111101100000000100",
    800 => "11011111111110111001111011111111",
    801 => "01100011111011111010110011100011",
    802 => "01111101110101100001001010001101",
    803 => "10101111111111110110000111011110",
    804 => "00111111110011110101000010100011",
    805 => "01110110011111100111010111100101",
    806 => "11110101110011100111010110100110",
    807 => "11101111111111101010100001111010",
    808 => "11101111111011101010010010110100",
    809 => "10111111110110111111100100011010",
    810 => "01111110101101110100001111110001",
    811 => "01011110100011110111111011010110",
    812 => "11011101001011111100111110100010",
    813 => "00100111111011100100010101000010",
    814 => "01111000010111110100010101110010",
    815 => "01111111011100011100101101100100",
    816 => "11111000110001110001111100010001",
    817 => "10111011111111111000010110111010",
    818 => "01101111101110110001010100001101",
    819 => "01111011110011101000001001100110",
    820 => "01111100011011000000011111110110",
    821 => "01110100111101111110011111001111",
    822 => "00001101111010110110011101110011",
    823 => "11101010110111011111100001010111",
    824 => "10111100010111011100011111011110",
    825 => "11101111111111011110111100010010",
    826 => "00111111101111011101011001001011",
    827 => "11011011100011011001011111011100",
    828 => "01111101111011110110011001011011",
    829 => "11111011101111111111001111100100",
    830 => "10111110111101111100000110111111",
    831 => "11000111011111011010101000000111",
    832 => "00101011111111110010111100010010",
    833 => "00110101011111110010010011000101",
    834 => "10111111111110110111010010101111",
    835 => "11111110011111101010100110000101",
    836 => "10110001111111111101110100101100",
    837 => "00110000111001100111000110000101",
    838 => "11110011101110000001000111001100",
    839 => "01101110111101111111011110010101",
    840 => "01100101111111110000001110100101",
    841 => "01110111111010110110110010111111",
    842 => "11100001111111100000101001111111",
    843 => "11001111101110100111010111110111",
    844 => "00100101001010110010000010000010",
    845 => "11001111111011111111000011000001",
    846 => "11111111011110010101011010000011",
    847 => "11100011000011010111001000000011",
    848 => "11001111111011111100000111101111",
    849 => "01111110111110010001000100000001",
    850 => "01010010111011100010010010110011",
    851 => "10111111011111110101101111010001",
    852 => "11010111111001111110001100011110",
    853 => "11011110011110110001111010010110",
    854 => "10111010111110111110001011010111",
    855 => "10111111011111010001100111000101",
    856 => "10101101110011010111111000010100",
    857 => "01111101010011111010000011100111",
    858 => "01110111111111100111001101010110",
    859 => "11101100001111111001100100010101",
    860 => "01101111111110100000011010110001",
    861 => "11111101111101101100100110001001",
    862 => "01001111011111001110111110100001",
    863 => "10110010101111101100011111100100",
    864 => "01111101110101110011011001101001",
    865 => "01010011011110111000001100101000",
    866 => "11100111110001110010001100010110",
    867 => "11111011111111101110010110100000",
    868 => "01001001011101110110100010110010",
    869 => "01110010110011010110001111101000",
    870 => "00011111101100110011000000111110",
    871 => "01111011001001011010000111110001",
    872 => "10111101010101111000101000101101",
    873 => "10111011011101111001001010001111",
    874 => "01111111010000110111100101011111",
    875 => "11011011111111000001001011011011",
    876 => "10010011011111010001000111110101",
    877 => "01011101111111111100111001100001",
    878 => "10011110111111100000001100011110",
    879 => "01001111111011101100011001110000",
    880 => "01111011110111111001011100000101",
    881 => "11111110111001111110110010001101",
    882 => "11110101101111110010101100110011",
    883 => "00101111000111110100010100011101",
    884 => "11110110010111110000110011001000",
    885 => "00111110111110111111001101001100",
    886 => "01111001111101111100010000000000",
    887 => "10111111111010101010000010111011",
    888 => "00111011111101110111001100111000",
    889 => "00101101011011011000000001001000",
    890 => "01111101111101100101111100000111",
    891 => "11110111011111110101001101110100",
    892 => "11101111111001010000111011111110",
    893 => "11111010001100010110011100011110",
    894 => "01101111001110111000000101000100",
    895 => "01011111111110001100100101001100",
    896 => "01011111011111100000100101100110",
    897 => "01111100111110100011110110001010",
    898 => "00100100111111011000010011001101",
    899 => "11001001110111010111101000101011",
    900 => "10111010111011100101111011101000",
    901 => "01111111001000001000011000101101",
    902 => "10010110011111101100111001111101",
    903 => "01110100110011110101011101001110",
    904 => "00111110011101010101010100011111",
    905 => "00101110100110110011110111000000",
    906 => "01101011110011111001001100001100",
    907 => "01111110111011111010100100111011",
    908 => "11111111011111110010010011111011",
    909 => "01111111010011111010011001100110",
    910 => "00111111111011011111000111000111",
    911 => "10111111111110011100010001011011",
    912 => "11101111111111101010110001111110",
    913 => "11111011001110111001000111110110",
    914 => "10111101111101110100000110010000",
    915 => "11011111111111011110010101001100",
    916 => "10111110110110110001111010011001",
    917 => "11110011101110011001010010011100",
    918 => "01111110010111111111001011101111",
    919 => "01001111101110110001110001001100",
    920 => "00111111011110010100111110010011",
    921 => "01111110111011111011100110000110",
    922 => "01011110111011111010100110000100",
    923 => "11011111111011110010001101001110",
    924 => "11110111101111111100110011001001",
    925 => "01111001011111101111111110110111",
    926 => "01111110001101110100010001100111",
    927 => "01111000101111111101101001001101",
    928 => "11101111110000111101001011011111",
    929 => "11010111011111110000101111010110",
    930 => "01110111011001111000010001100110",
    931 => "00110111110101010010010001111100",
    932 => "01111001000110110010110110111100",
    933 => "11111101111110110001011010111001",
    934 => "11111111010101011000101101110101",
    935 => "01011111100010101110111101100110",
    936 => "00111010111011101110001001011110",
    937 => "00101011111100101101001111010111",
    938 => "01110111001111111000011101101110",
    939 => "11110101101111111101101111001101",
    940 => "11010010101101111110010101011011",
    941 => "00111111101010011000011110111001",
    942 => "11011011110110000100100101001110",
    943 => "11011101011011100010101111101011",
    944 => "01111110111100110110111100000111",
    945 => "01011011111001110100011001000110",
    946 => "11110111100110100101001101010010",
    947 => "11111110110011110100110010011100",
    948 => "01111000001100011001010010101101",
    949 => "00011101001100111001110100010000",
    950 => "00111111111111010010110100000000",
    951 => "00111101111011110000101101010001",
    952 => "01110111110111100111111000010111",
    953 => "00011010110101110000100010100101",
    954 => "01101111101101011100001010100010",
    955 => "11001111010111111101101011110110",
    956 => "10100100110001001010110110101001",
    957 => "01011001100111101010010011110100",
    958 => "10010111111111110111100101101000",
    959 => "00111111111011101000100111100110",
    960 => "01011111001110101010011101111111",
    961 => "01110111000110110011001110110000",
    962 => "01111100110111010100011101000011",
    963 => "01100101111111011100110000101100",
    964 => "11111001111101110110001111000011",
    965 => "11101111110111100000011000110111",
    966 => "01100101010011110010110111011111",
    967 => "10110111100001010101011000110011",
    968 => "10011100110111010000111010100001",
    969 => "01101101110111110010010010000100",
    970 => "01110011111111110110001100110001",
    971 => "10111010001001100000110111011100",
    972 => "01011111010111011010101111000010",
    973 => "11110111111110010001110000100010",
    974 => "01000011111001110100011011110011",
    975 => "11111010111110110001001011100001",
    976 => "11011110111111111011011110111101",
    977 => "01000011111110110100001100000001",
    978 => "01101111111111110011111001111000",
    979 => "01100010101111110000001100101111",
    980 => "11011111111001110000100011100011",
    981 => "11110110110110110001000101010000",
    982 => "00111100011101110110110101000110",
    983 => "01110011110110111000000001011000",
    984 => "01100111111111111000010111101101",
    985 => "01110111111111110110001111111000",
    986 => "10001111111110101110101110110000",
    987 => "11110111111111110001101100001101",
    988 => "11111010000110110100010101100010",
    989 => "11011010010111111100101101110011",
    990 => "00011011001110101101110010100100",
    991 => "10111111101111011011001001101000",
    992 => "01111010111101010000011100011010",
    993 => "10001011010111111010111100010111",
    994 => "00111111111111101001001100011100",
    995 => "01100100011111010001001110110000",
    996 => "00101101111011011110111010111100",
    997 => "11011110001110100000101111101111",
    998 => "00101100010111110011110110111010",
    999 => "01110011111001111110110111001100");

  component fneg is
    port (A : in std_logic_vector (31 downto 0);
          CLK : in std_logic;
          Q : out std_logic_vector (31 downto 0));
  end component fneg;

  signal addr : integer :=  0;

  signal s_a : std_logic_vector (31 downto 0) := (others => '0');
  signal c : std_logic_vector (31 downto 0) := (others => '0');

  type buff is array (3 downto 0) of std_logic_vector (31 downto 0);
  signal cc : std_logic_vector (31 downto 0) := (others => '0');  
  signal QQ : std_logic_vector (7 downto 0) := x"2f";
  signal ccc : std_logic_vector (31 downto 0) := (others => '0'); 
  signal Q_buff : std_logic_vector (7 downto 0) := (others => '0');  
  signal state : std_logic_vector (1 downto 0) := (others => '0');
  signal i_isRunning : std_logic := 'U';
  signal i_result : std_logic := '1';
begin  -- architecture fneg_tb

  i_fneg : fneg port map (s_a,clk,c);
  isRunning <= i_isRunning;
  result <= i_result;

  ram_loop: process (clk,Q_buff) is
    variable ss : character;
    variable count : integer := 1;
  begin  -- process file_loop
    if clk'event and clk = '1' then    -- rising clock edge
      s_a <= a_lut (addr);
      cc <= ans_lut (addr);
      ccc <= cc ;

      if i_isRunning = '1' then  -- rising clock edge
        if ccc = c and i_result = '1' then
          i_result <= '1';
        else
          i_result <= '0';
        end if;
      end if;
      if addr >= array_max then
        if count > 0 then
          count := count - 1;
        else
          i_isRunning <= '0';
        end if;
      else
        if addr = 1 then
          i_isRunning <= '1';
        end if;
        addr <= addr + 1;
      end if;
    end if;

  end process ram_loop;

end architecture;
